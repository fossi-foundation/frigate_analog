magic
tech sky130A
magscale 1 2
timestamp 1719173892
<< checkpaint >>
rect 555256 92202 556228 92502
<< metal2 >>
rect 555256 92493 556228 92502
rect 555256 92211 555264 92493
rect 556219 92211 556228 92493
rect 555256 92202 556228 92211
<< via2 >>
rect 555264 92211 556219 92493
<< metal3 >>
rect 555256 92493 556228 92502
rect 555256 92211 555264 92493
rect 556219 92211 556228 92493
rect 555256 92202 556228 92211
<< end >>
