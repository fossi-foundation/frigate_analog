magic
tech sky130A
magscale 1 2
timestamp 1723648899
<< checkpaint >>
rect 70534 1051454 73254 1077338
rect 41200 1048875 81839 1051454
rect 39103 1039064 81839 1048875
rect 638072 1047955 986612 1185089
rect 637763 1047469 986612 1047955
rect 583513 1042008 624152 1043950
rect 583513 1039064 632284 1042008
rect 634122 1039064 986612 1047469
rect -1260 372718 986612 1039064
rect -1260 27767 719611 372718
rect -9140 -1260 719611 27767
rect -9140 -1876 630114 -1260
rect -384 -3036 630114 -1876
use analog_routes_bottom  analog_routes_bottom_0
timestamp 1717866854
transform 1 0 331431 0 1 40506
box 0 0 302118 22580
use analog_routes_left  analog_routes_left_0
timestamp 1723482278
transform 1 0 40451 0 1 349097
box 0 0 38119 501877
use analog_routes_right  analog_routes_right_0
timestamp 1722262877
transform 1 0 633291 0 1 50741
box 0 0 44160 800234
use analog_routes_top  analog_routes_top_0
timestamp 1717861592
transform 1 0 368282 0 1 966174
box 0 0 1800 30969
use analog_routes_user  analog_routes_user_0
timestamp 1723648899
transform 1 0 417670 0 1 830974
box 0 -20000 17024 20000
use analog_to_gpio_route  analog_to_gpio_route_0
timestamp 1717859832
transform 1 0 645945 0 1 863174
box 0 0 31376 2322
use analog_to_gpio_route  analog_to_gpio_route_1
timestamp 1717859832
transform -1 0 72020 0 1 879194
box 0 0 31376 2322
use analog_to_gpio_route  analog_to_gpio_route_2
timestamp 1717859832
transform -1 0 72020 0 1 900194
box 0 0 31376 2322
use analog_to_gpio_route  analog_to_gpio_route_3
timestamp 1717859832
transform -1 0 72020 0 1 921194
box 0 0 31376 2322
use analog_to_gpio_route  analog_to_gpio_route_4
timestamp 1717859832
transform -1 0 72020 0 1 942194
box 0 0 31376 2322
use analog_to_gpio_route  analog_to_gpio_route_5
timestamp 1717859832
transform 1 0 645945 0 1 926172
box 0 0 31376 2322
use analog_to_gpio_route  analog_to_gpio_route_6
timestamp 1717859832
transform 1 0 645945 0 1 905174
box 0 0 31376 2322
use analog_to_gpio_route  analog_to_gpio_route_7
timestamp 1717859832
transform 1 0 645945 0 1 884174
box 0 0 31376 2322
use analog_to_gpio_route_top  analog_to_gpio_route_top_0
timestamp 1717859897
transform 1 0 151882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_1
timestamp 1717859897
transform 1 0 79882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_2
timestamp 1717859897
transform 1 0 103882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_3
timestamp 1717859897
transform 1 0 127882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_4
timestamp 1717859897
transform 1 0 245882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_5
timestamp 1717859897
transform 1 0 221882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_6
timestamp 1717859897
transform 1 0 293882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_7
timestamp 1717859897
transform 1 0 269882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_8
timestamp 1717859897
transform 1 0 359882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_9
timestamp 1717859897
transform 1 0 336882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_10
timestamp 1717859897
transform 1 0 456882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_11
timestamp 1717859897
transform 1 0 432882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_12
timestamp 1717859897
transform 1 0 504882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_13
timestamp 1717859897
transform 1 0 480882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_14
timestamp 1717859897
transform 1 0 574882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_16
timestamp 1717859897
transform 1 0 598882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_route_top  analog_to_gpio_route_top_17
timestamp 1717859897
transform 1 0 622882 0 1 966174
box 0 0 1401 31117
use analog_to_gpio_top_right  analog_to_gpio_top_right_0
timestamp 1723482457
transform 1 0 640770 0 1 966174
box -6 0 7162 31606
use frigate_analog  frigate_analog_0
timestamp 1723485911
transform 1 0 71670 0 1 850974
box -6 -20 574622 115224
use frigate_timing_frontend  frigate_timing_frontend_0
timestamp 1719949696
transform 1 0 247240 0 1 41166
box 1 -21 84200 25600
use panamax  panamax_0 ../dependencies/panamax/mag
timestamp 1719158962
transform 1 0 151 0 1 204
box -151 -204 717751 1037600
<< end >>
