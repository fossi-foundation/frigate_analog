magic
tech sky130A
magscale 1 2
timestamp 1724602578
<< checkpaint >>
rect -1302 33010 1906 33364
rect -1702 31680 8720 33010
rect -1702 30838 8772 31680
rect -1702 28320 9044 30838
rect -1260 -1260 2661 28320
rect 4284 28126 9044 28320
rect 4852 -1260 8773 28126
rect -642030 -967434 -639509 -964913
<< metal2 >>
rect 6742 31091 7056 31117
rect 6742 30712 6775 31091
rect 7024 30712 7056 31091
rect 6742 30683 7056 30712
<< via2 >>
rect 6775 30712 7024 31091
<< metal3 >>
rect 6712 31091 7162 31117
rect 6712 30932 6775 31091
rect 7024 30932 7162 31091
rect 6712 30642 6740 30932
rect 7134 30642 7162 30932
<< via3 >>
rect 6740 30712 6775 30932
rect 6775 30712 7024 30932
rect 7024 30712 7134 30932
rect 6740 30516 7134 30712
<< metal4 >>
rect 0 949 200 31448
rect 6712 30932 7162 30957
rect 0 905 320 949
rect 0 194 38 905
rect 279 194 320 905
rect 0 149 320 194
rect 600 0 800 30766
rect 6712 30516 6740 30932
rect 7134 30516 7162 30932
rect 6712 30482 7162 30516
rect 1200 949 1400 30050
rect 1080 903 1400 949
rect 1080 192 1121 903
rect 1362 192 1400 903
rect 1080 149 1400 192
<< via4 >>
rect 38 194 279 905
rect 1121 192 1362 903
<< metal5 >>
rect 0 31268 7160 31588
rect 600 30562 7162 30882
rect 1200 29868 7160 30188
rect 0 905 1401 949
rect 0 194 38 905
rect 279 903 1401 905
rect 279 194 1121 903
rect 0 192 1121 194
rect 1362 192 1401 903
rect 0 149 1401 192
use cv3_via4_2cut  cv3_via4_2cut_0
timestamp 1717863568
transform 1 0 6470 0 1 30564
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_1
timestamp 1717863568
transform 1 0 -6 0 1 31238
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_2
timestamp 1717863568
transform 1 0 600 0 1 30528
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_3
timestamp 1717863568
transform 1 0 1196 0 1 29830
box 0 0 688 368
<< properties >>
string FIXED_BBOX 0 0 7162 31588
string LEFclass COVER
<< end >>
