magic
tech sky130A
magscale 1 2
timestamp 1724444698
<< metal1 >>
rect -41 13354 122 13375
rect -41 13004 -25 13354
rect 107 13004 122 13354
rect 885 13356 1048 13374
rect 885 13006 902 13356
rect 1034 13006 1048 13356
rect 885 13005 1048 13006
rect 4581 13354 4745 13369
rect -41 12989 122 13004
rect 4581 13004 4601 13354
rect 4733 13004 4745 13354
rect 5513 13356 5677 13367
rect 5513 13006 5528 13356
rect 5660 13006 5677 13356
rect 5513 13004 5677 13006
rect 9207 13354 9371 13367
rect 9207 13004 9227 13354
rect 9359 13004 9371 13354
rect 4581 13002 4745 13004
rect 9207 13002 9371 13004
rect 10139 13356 10303 13367
rect 10139 13006 10154 13356
rect 10286 13271 10303 13356
rect 13833 13354 13997 13367
rect 10286 13009 10305 13271
rect 10286 13006 10303 13009
rect 10139 13002 10303 13006
rect 13833 13004 13853 13354
rect 13985 13004 13997 13354
rect 14765 13356 14929 13367
rect 14765 13006 14780 13356
rect 14912 13271 14929 13356
rect 18459 13354 18623 13367
rect 14912 13009 14931 13271
rect 18459 13260 18479 13354
rect 14912 13006 14929 13009
rect 14765 13004 14929 13006
rect 18457 13004 18479 13260
rect 18611 13004 18623 13354
rect 13833 13002 13997 13004
rect 18457 12989 18623 13004
rect 19391 13356 19555 13367
rect 19391 13006 19406 13356
rect 19538 13271 19555 13356
rect 23085 13354 23249 13367
rect 19538 13009 19557 13271
rect 19538 13006 19555 13009
rect 18457 12987 18608 12989
rect 19391 12987 19555 13006
rect 23085 13004 23105 13354
rect 23237 13004 23249 13354
rect 24017 13356 24181 13367
rect 24017 13006 24032 13356
rect 24164 13271 24181 13356
rect 27711 13354 27875 13367
rect 24164 13009 24183 13271
rect 24164 13006 24181 13009
rect 24017 13005 24181 13006
rect 23085 13002 23249 13004
rect 27711 13004 27731 13354
rect 27863 13004 27875 13354
rect 27711 13003 27875 13004
rect 28643 13356 28807 13367
rect 28643 13006 28658 13356
rect 28790 13271 28807 13356
rect 32337 13354 32501 13367
rect 28790 13009 28809 13271
rect 28790 13006 28807 13009
rect 28643 13002 28807 13006
rect 32337 13004 32357 13354
rect 32489 13004 32501 13354
rect 32337 13003 32501 13004
rect 33269 13356 33433 13367
rect 33269 13006 33284 13356
rect 33416 13271 33433 13356
rect 36963 13354 37127 13367
rect 33416 13009 33435 13271
rect 33416 13006 33433 13009
rect 33269 13003 33433 13006
rect 36963 13004 36983 13354
rect 37115 13004 37127 13354
rect 37895 13356 38059 13367
rect 37895 13006 37910 13356
rect 38042 13271 38059 13356
rect 41589 13354 41753 13367
rect 41589 13293 41609 13354
rect 38042 13009 38061 13271
rect 38042 13006 38059 13009
rect 37895 13005 38059 13006
rect 36963 13003 37127 13004
rect 41587 13004 41609 13293
rect 41741 13004 41753 13354
rect 41587 12989 41753 13004
rect 42521 13356 42685 13367
rect 42521 13006 42536 13356
rect 42668 13271 42685 13356
rect 46215 13354 46379 13367
rect 42668 13009 42687 13271
rect 42668 13006 42685 13009
rect 41587 12987 41738 12989
rect 42521 12987 42685 13006
rect 46215 13004 46235 13354
rect 46367 13004 46379 13354
rect 47147 13356 47311 13367
rect 47147 13006 47162 13356
rect 47294 13271 47311 13356
rect 50841 13354 51005 13367
rect 47294 13009 47313 13271
rect 47294 13006 47311 13009
rect 47147 13004 47311 13006
rect 50841 13004 50861 13354
rect 50993 13004 51005 13354
rect 51773 13356 51937 13367
rect 51773 13006 51788 13356
rect 51920 13271 51937 13356
rect 55467 13354 55631 13367
rect 51920 13009 51939 13271
rect 51920 13006 51937 13009
rect 51773 13005 51937 13006
rect 46215 13003 46379 13004
rect 50841 13003 51005 13004
rect 55467 13004 55487 13354
rect 55619 13004 55631 13354
rect 55467 13003 55631 13004
rect 56399 13356 56563 13367
rect 56399 13006 56414 13356
rect 56546 13271 56563 13356
rect 60093 13354 60257 13367
rect 56546 13009 56565 13271
rect 56546 13006 56563 13009
rect 56399 13003 56563 13006
rect 60093 13004 60113 13354
rect 60245 13004 60257 13354
rect 61025 13356 61189 13367
rect 61025 13006 61040 13356
rect 61172 13271 61189 13356
rect 64719 13354 64883 13367
rect 64719 13285 64739 13354
rect 61172 13009 61191 13271
rect 61172 13006 61189 13009
rect 61025 13004 61189 13006
rect 64717 13004 64739 13285
rect 64871 13004 64883 13354
rect 60093 13002 60257 13004
rect 64717 12989 64883 13004
rect 65651 13356 65815 13367
rect 65651 13006 65666 13356
rect 65798 13271 65815 13356
rect 69345 13354 69509 13367
rect 65798 13009 65817 13271
rect 65798 13006 65815 13009
rect 64717 12987 64868 12989
rect 65651 12987 65815 13006
rect 69345 13004 69365 13354
rect 69497 13004 69509 13354
rect 69345 13002 69509 13004
rect 70277 13356 70441 13367
rect 70277 13006 70292 13356
rect 70424 13271 70441 13356
rect 73971 13354 74135 13367
rect 70424 13009 70443 13271
rect 70424 13006 70441 13009
rect 70277 13003 70441 13006
rect 73971 13004 73991 13354
rect 74123 13004 74135 13354
rect 74903 13356 75067 13367
rect 74903 13006 74918 13356
rect 75050 13271 75067 13356
rect 78597 13354 78761 13367
rect 75050 13009 75069 13271
rect 75050 13006 75067 13009
rect 74903 13004 75067 13006
rect 78597 13004 78617 13354
rect 78749 13004 78761 13354
rect 79529 13356 79693 13367
rect 79529 13006 79544 13356
rect 79676 13271 79693 13356
rect 83223 13354 83387 13367
rect 79676 13009 79695 13271
rect 79676 13006 79693 13009
rect 79529 13004 79693 13006
rect 83223 13004 83243 13354
rect 83375 13004 83387 13354
rect 73971 13002 74135 13004
rect 78597 13002 78761 13004
rect 83223 13002 83387 13004
rect 84155 13356 84319 13367
rect 84155 13006 84170 13356
rect 84302 13271 84319 13356
rect 87849 13354 88013 13367
rect 87849 13285 87869 13354
rect 84302 13009 84321 13271
rect 84302 13006 84319 13009
rect 84155 13003 84319 13006
rect 87847 13004 87869 13285
rect 88001 13004 88013 13354
rect 87847 12989 88013 13004
rect 88781 13356 88945 13367
rect 88781 13006 88796 13356
rect 88928 13271 88945 13356
rect 92475 13354 92639 13367
rect 88928 13009 88947 13271
rect 88928 13006 88945 13009
rect 87847 12987 87998 12989
rect 88781 12987 88945 13006
rect 92475 13004 92495 13354
rect 92627 13004 92639 13354
rect 93407 13356 93571 13367
rect 93407 13006 93422 13356
rect 93554 13271 93571 13356
rect 97101 13354 97265 13367
rect 93554 13009 93573 13271
rect 93554 13006 93571 13009
rect 93407 13004 93571 13006
rect 97101 13004 97121 13354
rect 97253 13004 97265 13354
rect 98033 13356 98197 13367
rect 98033 13006 98048 13356
rect 98180 13271 98197 13356
rect 101727 13354 101891 13367
rect 98180 13009 98199 13271
rect 98180 13006 98197 13009
rect 98033 13004 98197 13006
rect 101727 13004 101747 13354
rect 101879 13004 101891 13354
rect 102659 13356 102823 13367
rect 102659 13006 102674 13356
rect 102806 13271 102823 13356
rect 106353 13354 106517 13367
rect 106353 13317 106373 13354
rect 102806 13009 102825 13271
rect 102806 13006 102823 13009
rect 102659 13005 102823 13006
rect 92475 13003 92639 13004
rect 97101 13003 97265 13004
rect 101727 13002 101891 13004
rect 106351 13004 106373 13317
rect 106505 13004 106517 13354
rect 106351 12989 106517 13004
rect 107285 13356 107449 13367
rect 107285 13006 107300 13356
rect 107432 13271 107449 13356
rect 110979 13354 111143 13367
rect 107432 13009 107451 13271
rect 107432 13006 107449 13009
rect 106351 12987 106502 12989
rect 107285 12987 107449 13006
rect 110979 13004 110999 13354
rect 111131 13004 111143 13354
rect 111911 13356 112075 13367
rect 111911 13006 111926 13356
rect 112058 13271 112075 13356
rect 115605 13354 115769 13367
rect 112058 13009 112077 13271
rect 112058 13006 112075 13009
rect 111911 13004 112075 13006
rect 115605 13004 115625 13354
rect 115757 13004 115769 13354
rect 116537 13356 116701 13367
rect 116537 13006 116552 13356
rect 116684 13271 116701 13356
rect 120231 13354 120395 13367
rect 116684 13009 116703 13271
rect 120231 13252 120251 13354
rect 116684 13006 116701 13009
rect 116537 13004 116701 13006
rect 120229 13004 120251 13252
rect 120383 13004 120395 13354
rect 110979 13003 111143 13004
rect 115605 13003 115769 13004
rect 120229 12989 120395 13004
rect 121163 13356 121327 13367
rect 121163 13006 121178 13356
rect 121310 13271 121327 13356
rect 124857 13354 125021 13367
rect 121310 13009 121329 13271
rect 121310 13006 121327 13009
rect 120229 12987 120380 12989
rect 121163 12987 121327 13006
rect 124857 13004 124877 13354
rect 125009 13004 125021 13354
rect 125789 13356 125953 13367
rect 125789 13006 125804 13356
rect 125936 13271 125953 13356
rect 129483 13354 129647 13367
rect 125936 13009 125955 13271
rect 125936 13006 125953 13009
rect 125789 13004 125953 13006
rect 129483 13004 129503 13354
rect 129635 13004 129647 13354
rect 130415 13356 130579 13367
rect 130415 13006 130430 13356
rect 130562 13271 130579 13356
rect 134109 13314 134273 13327
rect 130562 13009 130581 13271
rect 134109 13245 134129 13314
rect 130562 13006 130579 13009
rect 130415 13004 130579 13006
rect 124857 13002 125021 13004
rect 129483 13002 129647 13004
rect -47 7457 101 9928
rect 945 7503 1002 10753
rect 4579 7471 4727 9977
rect 5571 7546 5628 10764
rect 9205 7471 9353 9944
rect 10197 7519 10254 10796
rect 13831 7440 13979 9923
rect 14823 7552 14880 10796
rect 18457 7458 18605 12987
rect 19446 7503 19554 12987
rect 23083 7471 23231 9901
rect 24075 7465 24132 10780
rect 27709 7471 27857 9961
rect 28701 7503 28758 10796
rect 32335 7446 32483 9950
rect 33327 7552 33384 10775
rect 36961 7457 37109 9961
rect 37953 7492 38010 10764
rect 41587 7471 41735 12987
rect 42576 7487 42684 12987
rect 46213 7471 46361 9972
rect 47205 7535 47262 10780
rect 50839 7471 50987 9972
rect 51831 7524 51888 10764
rect 55465 7467 55613 9950
rect 56457 7486 56514 10769
rect 60091 7451 60239 10059
rect 61083 7546 61140 10775
rect 64717 7471 64865 12987
rect 65706 7487 65814 12987
rect 69343 7471 69491 9928
rect 70335 7519 70392 10747
rect 73969 7471 74117 9923
rect 74961 7541 75018 10764
rect 78595 7457 78743 9917
rect 79587 7590 79644 10740
rect 83221 7471 83369 9944
rect 84213 7524 84270 10747
rect 87847 7471 87995 12987
rect 88836 7470 88944 12987
rect 92473 7471 92621 9966
rect 93465 7519 93522 10769
rect 97099 7471 97247 9966
rect 98091 7497 98148 10758
rect 101725 7471 101873 9944
rect 102717 7541 102774 10769
rect 106351 7458 106499 12987
rect 107340 7478 107448 12987
rect 110977 7471 111125 10037
rect 111969 7470 112026 10769
rect 115603 7435 115751 9977
rect 116595 7497 116652 10758
rect 120229 7450 120377 12987
rect 121218 7510 121326 12987
rect 134107 12964 134129 13245
rect 134261 12964 134273 13314
rect 134107 12949 134273 12964
rect 135041 13316 135205 13327
rect 135041 12966 135056 13316
rect 135188 13231 135205 13316
rect 135188 12969 135207 13231
rect 135188 12966 135205 12969
rect 134107 12947 134258 12949
rect 135041 12947 135205 12966
rect 124855 7471 125003 9928
rect 125847 7475 125904 10769
rect 129481 7471 129629 9939
rect 130473 7513 130530 10769
rect 134107 7471 134255 12947
rect 135096 7487 135204 12947
<< via1 >>
rect -25 13004 107 13354
rect 902 13006 1034 13356
rect 4601 13004 4733 13354
rect 5528 13006 5660 13356
rect 9227 13004 9359 13354
rect 10154 13006 10286 13356
rect 13853 13004 13985 13354
rect 14780 13006 14912 13356
rect 18479 13004 18611 13354
rect 19406 13006 19538 13356
rect 23105 13004 23237 13354
rect 24032 13006 24164 13356
rect 27731 13004 27863 13354
rect 28658 13006 28790 13356
rect 32357 13004 32489 13354
rect 33284 13006 33416 13356
rect 36983 13004 37115 13354
rect 37910 13006 38042 13356
rect 41609 13004 41741 13354
rect 42536 13006 42668 13356
rect 46235 13004 46367 13354
rect 47162 13006 47294 13356
rect 50861 13004 50993 13354
rect 51788 13006 51920 13356
rect 55487 13004 55619 13354
rect 56414 13006 56546 13356
rect 60113 13004 60245 13354
rect 61040 13006 61172 13356
rect 64739 13004 64871 13354
rect 65666 13006 65798 13356
rect 69365 13004 69497 13354
rect 70292 13006 70424 13356
rect 73991 13004 74123 13354
rect 74918 13006 75050 13356
rect 78617 13004 78749 13354
rect 79544 13006 79676 13356
rect 83243 13004 83375 13354
rect 84170 13006 84302 13356
rect 87869 13004 88001 13354
rect 88796 13006 88928 13356
rect 92495 13004 92627 13354
rect 93422 13006 93554 13356
rect 97121 13004 97253 13354
rect 98048 13006 98180 13356
rect 101747 13004 101879 13354
rect 102674 13006 102806 13356
rect 106373 13004 106505 13354
rect 107300 13006 107432 13356
rect 110999 13004 111131 13354
rect 111926 13006 112058 13356
rect 115625 13004 115757 13354
rect 116552 13006 116684 13356
rect 120251 13004 120383 13354
rect 121178 13006 121310 13356
rect 124877 13004 125009 13354
rect 125804 13006 125936 13356
rect 129503 13004 129635 13354
rect 130430 13006 130562 13356
rect 134129 12964 134261 13314
rect 135056 12966 135188 13316
<< metal2 >>
rect 25403 16286 25593 16287
rect 28641 16286 28806 16287
rect -215 16247 122 16282
rect -215 15940 -183 16247
rect 88 15940 122 16247
rect -215 15912 122 15940
rect 881 16259 1218 16286
rect 881 15952 910 16259
rect 1181 15952 1218 16259
rect 881 15916 1218 15952
rect 2129 16263 2466 16286
rect 2129 15956 2161 16263
rect 2432 15956 2466 16263
rect 2129 15916 2466 15956
rect 3753 16255 4090 16286
rect 3753 15948 3784 16255
rect 4055 15948 4090 16255
rect 3753 15916 4090 15948
rect 4411 16247 4748 16282
rect 4411 15940 4443 16247
rect 4714 15940 4748 16247
rect -44 13354 120 15912
rect -44 13004 -25 13354
rect 107 13004 120 13354
rect -44 12989 120 13004
rect 885 13356 1050 15916
rect 885 13006 902 13356
rect 1034 13006 1050 13356
rect 2273 13086 2463 15916
rect 885 12988 1050 13006
rect 2608 11630 3040 13889
rect 3755 13104 3923 15916
rect 4411 15912 4748 15940
rect 5507 16259 5844 16286
rect 5507 15952 5536 16259
rect 5807 15952 5844 16259
rect 5507 15916 5844 15952
rect 6755 16263 7092 16286
rect 6755 15956 6787 16263
rect 7058 15956 7092 16263
rect 6755 15916 7092 15956
rect 8379 16255 8716 16286
rect 8379 15948 8410 16255
rect 8681 15948 8716 16255
rect 8379 15916 8716 15948
rect 9037 16247 9374 16282
rect 9037 15940 9069 16247
rect 9340 15940 9374 16247
rect 4582 13354 4746 15912
rect 4582 13004 4601 13354
rect 4733 13004 4746 13354
rect 4582 12989 4746 13004
rect 5511 13356 5676 15916
rect 5511 13006 5528 13356
rect 5660 13006 5676 13356
rect 5511 12988 5676 13006
rect 6899 12982 7089 15916
rect 8381 12962 8549 15916
rect 9037 15912 9374 15940
rect 10133 16259 10470 16286
rect 10133 15952 10162 16259
rect 10433 15952 10470 16259
rect 10133 15916 10470 15952
rect 11381 16263 11718 16286
rect 11381 15956 11413 16263
rect 11684 15956 11718 16263
rect 11381 15916 11718 15956
rect 13005 16255 13342 16286
rect 13863 16281 14200 16282
rect 13005 15948 13036 16255
rect 13307 15948 13342 16255
rect 13005 15916 13342 15948
rect 13834 16247 14200 16281
rect 13834 15940 13895 16247
rect 14166 15940 14200 16247
rect 9208 13354 9372 15912
rect 9208 13004 9227 13354
rect 9359 13004 9372 13354
rect 9208 12989 9372 13004
rect 10137 13356 10302 15916
rect 10137 13006 10154 13356
rect 10286 13006 10302 13356
rect 10137 12988 10302 13006
rect 11525 12982 11715 15916
rect 13007 12962 13175 15916
rect 13834 15912 14200 15940
rect 14759 16259 15096 16286
rect 14759 15952 14788 16259
rect 15059 15952 15096 16259
rect 14759 15916 15096 15952
rect 16007 16263 16344 16286
rect 16007 15956 16039 16263
rect 16310 15956 16344 16263
rect 16007 15916 16344 15956
rect 17631 16255 17968 16286
rect 17631 15948 17662 16255
rect 17933 15948 17968 16255
rect 17631 15916 17968 15948
rect 18289 16247 18626 16282
rect 18289 15940 18321 16247
rect 18592 15940 18626 16247
rect 13834 13354 13998 15912
rect 13834 13004 13853 13354
rect 13985 13004 13998 13354
rect 13834 12989 13998 13004
rect 14763 13356 14928 15916
rect 14763 13006 14780 13356
rect 14912 13006 14928 13356
rect 14763 12988 14928 13006
rect 16151 12982 16341 15916
rect 17633 12962 17801 15916
rect 18289 15912 18626 15940
rect 19385 16259 19722 16286
rect 19385 15952 19414 16259
rect 19685 15952 19722 16259
rect 19385 15916 19722 15952
rect 20633 16263 20970 16286
rect 20633 15956 20665 16263
rect 20936 15956 20970 16263
rect 20633 15916 20970 15956
rect 22257 16255 22594 16286
rect 22257 15948 22288 16255
rect 22559 15948 22594 16255
rect 22257 15916 22594 15948
rect 22915 16247 23252 16282
rect 22915 15940 22947 16247
rect 23218 15940 23252 16247
rect 18460 13354 18624 15912
rect 18460 13004 18479 13354
rect 18611 13004 18624 13354
rect 18460 12989 18624 13004
rect 19389 13356 19554 15916
rect 19389 13006 19406 13356
rect 19538 13006 19554 13356
rect 20777 13265 20967 15916
rect 22259 13287 22427 15916
rect 22915 15912 23252 15940
rect 24011 16259 24348 16286
rect 24011 15952 24040 16259
rect 24311 15952 24348 16259
rect 24011 15916 24348 15952
rect 25403 16263 25906 16286
rect 25403 15956 25601 16263
rect 25872 15956 25906 16263
rect 25403 15916 25906 15956
rect 26283 16255 26620 16286
rect 26283 15948 26314 16255
rect 26585 16081 26620 16255
rect 27481 16247 27876 16282
rect 26585 15948 27053 16081
rect 26283 15916 27053 15948
rect 19389 12988 19554 13006
rect 20774 12982 20967 13265
rect 2270 7433 2460 9876
rect 3168 434 3600 12133
rect 3752 7451 3920 9859
rect 6896 7433 7086 9903
rect 7794 412 8226 12133
rect 11860 11723 12292 12786
rect 8378 7451 8546 9881
rect 11522 7433 11712 9892
rect 12420 432 12852 12133
rect 13004 7451 13172 9902
rect 16148 7433 16338 9870
rect 16486 7206 16918 8764
rect 17046 494 17478 12133
rect 17630 7451 17798 9854
rect 20774 7433 20964 12982
rect 22256 12962 22427 13287
rect 23086 13354 23250 15912
rect 23086 13004 23105 13354
rect 23237 13004 23250 13354
rect 23086 12989 23250 13004
rect 24015 13356 24180 15916
rect 24015 13006 24032 13356
rect 24164 13006 24180 13356
rect 24015 12988 24180 13006
rect 25403 12982 25593 15916
rect 21112 7167 21544 10816
rect 22256 7451 22424 12962
rect 25741 12793 26173 13287
rect 26885 12962 27053 15916
rect 27481 15940 27513 16247
rect 27784 15940 27876 16247
rect 27481 15912 27876 15940
rect 27712 13354 27876 15912
rect 27712 13004 27731 13354
rect 27863 13004 27876 13354
rect 27712 12989 27876 13004
rect 28641 16259 29074 16286
rect 28641 15952 28766 16259
rect 29037 15952 29074 16259
rect 28641 15916 29074 15952
rect 29885 16263 30222 16286
rect 29885 15956 29917 16263
rect 30188 15956 30222 16263
rect 29885 15916 30222 15956
rect 31509 16255 31846 16286
rect 31509 15948 31540 16255
rect 31811 15948 31846 16255
rect 31509 15916 31846 15948
rect 32167 16247 32504 16282
rect 32167 15940 32199 16247
rect 32470 15940 32504 16247
rect 28641 13356 28806 15916
rect 28641 13006 28658 13356
rect 28790 13006 28806 13356
rect 28641 12988 28806 13006
rect 30029 12982 30219 15916
rect 31511 12962 31679 15916
rect 32167 15912 32504 15940
rect 33263 16259 33600 16286
rect 33263 15952 33292 16259
rect 33563 15952 33600 16259
rect 33263 15916 33600 15952
rect 34511 16263 34848 16286
rect 34511 15956 34543 16263
rect 34814 15956 34848 16263
rect 34511 15916 34848 15956
rect 36135 16255 36472 16286
rect 36135 15948 36166 16255
rect 36437 15948 36472 16255
rect 36135 15916 36472 15948
rect 36793 16247 37130 16282
rect 36793 15940 36825 16247
rect 37096 15940 37130 16247
rect 32338 13354 32502 15912
rect 32338 13004 32357 13354
rect 32489 13004 32502 13354
rect 32338 12989 32502 13004
rect 33267 13356 33432 15916
rect 33267 13006 33284 13356
rect 33416 13006 33432 13356
rect 33267 12988 33432 13006
rect 34655 12982 34845 15916
rect 36137 12962 36305 15916
rect 36793 15912 37130 15940
rect 37889 16259 38226 16286
rect 37889 15952 37918 16259
rect 38189 15952 38226 16259
rect 37889 15916 38226 15952
rect 39137 16263 39474 16286
rect 39137 15956 39169 16263
rect 39440 15956 39474 16263
rect 39137 15916 39474 15956
rect 40761 16255 41098 16286
rect 40761 15948 40792 16255
rect 41063 15948 41098 16255
rect 40761 15916 41098 15948
rect 41419 16247 41756 16282
rect 41419 15940 41451 16247
rect 41722 15940 41756 16247
rect 36964 13354 37128 15912
rect 36964 13004 36983 13354
rect 37115 13004 37128 13354
rect 36964 12989 37128 13004
rect 37893 13356 38058 15916
rect 37893 13006 37910 13356
rect 38042 13006 38058 13356
rect 37893 12988 38058 13006
rect 39281 12982 39471 15916
rect 40763 12962 40931 15916
rect 41419 15912 41756 15940
rect 42515 16259 42852 16286
rect 42515 15952 42544 16259
rect 42815 15952 42852 16259
rect 42515 15916 42852 15952
rect 43763 16263 44100 16286
rect 43763 15956 43795 16263
rect 44066 15956 44100 16263
rect 43763 15916 44100 15956
rect 45387 16255 45724 16286
rect 45387 15948 45418 16255
rect 45689 15948 45724 16255
rect 45387 15916 45724 15948
rect 46045 16247 46382 16282
rect 46045 15940 46077 16247
rect 46348 15940 46382 16247
rect 41590 13354 41754 15912
rect 41590 13004 41609 13354
rect 41741 13004 41754 13354
rect 41590 12989 41754 13004
rect 42519 13356 42684 15916
rect 42519 13006 42536 13356
rect 42668 13006 42684 13356
rect 43907 13289 44097 15916
rect 42519 12988 42684 13006
rect 43904 12982 44097 13289
rect 45389 13287 45557 15916
rect 46045 15912 46382 15940
rect 47141 16259 47478 16286
rect 47141 15952 47170 16259
rect 47441 15952 47478 16259
rect 47141 15916 47478 15952
rect 48389 16263 48726 16286
rect 48389 15956 48421 16263
rect 48692 15956 48726 16263
rect 48389 15916 48726 15956
rect 50013 16255 50350 16286
rect 50013 15948 50044 16255
rect 50315 15948 50350 16255
rect 50013 15916 50350 15948
rect 50671 16247 51008 16282
rect 50671 15940 50703 16247
rect 50974 15940 51008 16247
rect 25400 7433 25590 9959
rect 21672 520 22104 7087
rect 26302 924 26734 12133
rect 26882 7451 27050 9937
rect 30026 7433 30216 9937
rect 30928 972 31360 12133
rect 31508 7425 31676 9904
rect 34652 7433 34842 9861
rect 35550 934 35982 12133
rect 36134 7446 36302 9872
rect 39278 7433 39468 9872
rect 39619 9157 40051 10210
rect 39616 7205 40048 8139
rect 40176 934 40608 12133
rect 40760 7451 40928 9904
rect 43904 7433 44094 12982
rect 45386 12962 45557 13287
rect 46216 13354 46380 15912
rect 46216 13004 46235 13354
rect 46367 13004 46380 13354
rect 46216 12989 46380 13004
rect 47145 13356 47310 15916
rect 47145 13006 47162 13356
rect 47294 13006 47310 13356
rect 47145 12988 47310 13006
rect 48533 12982 48723 15916
rect 44242 7195 44674 10178
rect 45386 7451 45554 12962
rect 48871 12825 49303 13843
rect 50015 12962 50183 15916
rect 50671 15912 51008 15940
rect 51767 16259 52104 16286
rect 51767 15952 51796 16259
rect 52067 15952 52104 16259
rect 51767 15916 52104 15952
rect 53015 16263 53352 16286
rect 53015 15956 53047 16263
rect 53318 15956 53352 16263
rect 53015 15916 53352 15956
rect 54639 16255 54976 16286
rect 54639 15948 54670 16255
rect 54941 15948 54976 16255
rect 54639 15916 54976 15948
rect 55297 16247 55634 16282
rect 55297 15940 55329 16247
rect 55600 15940 55634 16247
rect 50842 13354 51006 15912
rect 50842 13004 50861 13354
rect 50993 13004 51006 13354
rect 50842 12989 51006 13004
rect 51771 13356 51936 15916
rect 51771 13006 51788 13356
rect 51920 13006 51936 13356
rect 51771 12988 51936 13006
rect 53159 12982 53349 15916
rect 54641 12962 54809 15916
rect 55297 15912 55634 15940
rect 56393 16259 56730 16286
rect 56393 15952 56422 16259
rect 56693 15952 56730 16259
rect 56393 15916 56730 15952
rect 57641 16263 57978 16286
rect 57641 15956 57673 16263
rect 57944 15956 57978 16263
rect 57641 15916 57978 15956
rect 59265 16255 59602 16286
rect 59265 15948 59296 16255
rect 59567 15948 59602 16255
rect 59265 15916 59602 15948
rect 59923 16247 60260 16282
rect 59923 15940 59955 16247
rect 60226 15940 60260 16247
rect 55468 13354 55632 15912
rect 55468 13004 55487 13354
rect 55619 13004 55632 13354
rect 55468 12989 55632 13004
rect 56397 13356 56562 15916
rect 56397 13006 56414 13356
rect 56546 13006 56562 13356
rect 56397 12988 56562 13006
rect 57785 12982 57975 15916
rect 59267 12962 59435 15916
rect 59923 15912 60260 15940
rect 61019 16259 61356 16286
rect 61019 15952 61048 16259
rect 61319 15952 61356 16259
rect 61019 15916 61356 15952
rect 61867 16263 62204 16286
rect 61867 15956 61899 16263
rect 62170 16093 62204 16263
rect 64191 16255 64528 16286
rect 64191 16096 64222 16255
rect 62170 15956 62602 16093
rect 61867 15916 62602 15956
rect 63893 15948 64222 16096
rect 64493 15948 64528 16255
rect 63893 15916 64528 15948
rect 64720 16247 65186 16282
rect 64720 15940 64881 16247
rect 65152 15940 65186 16247
rect 60094 13354 60258 15912
rect 60094 13004 60113 13354
rect 60245 13004 60258 13354
rect 60094 12989 60258 13004
rect 61023 13356 61188 15916
rect 61023 13006 61040 13356
rect 61172 13006 61188 13356
rect 61023 12988 61188 13006
rect 62411 12982 62601 15916
rect 63893 12962 64061 15916
rect 64720 15912 65186 15940
rect 65645 16259 65982 16286
rect 65645 15952 65674 16259
rect 65945 15952 65982 16259
rect 65645 15916 65982 15952
rect 67037 16263 67411 16286
rect 67037 15956 67106 16263
rect 67377 15956 67411 16263
rect 67037 15916 67411 15956
rect 68517 16255 68854 16286
rect 68517 15948 68548 16255
rect 68819 15948 68854 16255
rect 68517 15916 68854 15948
rect 69175 16247 69512 16282
rect 69175 15940 69207 16247
rect 69478 15940 69512 16247
rect 64720 13354 64884 15912
rect 64720 13004 64739 13354
rect 64871 13004 64884 13354
rect 64720 12989 64884 13004
rect 65649 13356 65814 15916
rect 65649 13006 65666 13356
rect 65798 13006 65814 13356
rect 67037 13265 67227 15916
rect 68519 13303 68687 15916
rect 69175 15912 69512 15940
rect 70271 16259 70608 16286
rect 70271 15952 70300 16259
rect 70571 15952 70608 16259
rect 70271 15916 70608 15952
rect 71519 16263 71856 16286
rect 71519 15956 71551 16263
rect 71822 15956 71856 16263
rect 71519 15916 71856 15956
rect 73143 16255 73480 16286
rect 73143 15948 73174 16255
rect 73445 15948 73480 16255
rect 73143 15916 73480 15948
rect 73971 16247 74308 16282
rect 73971 15940 74003 16247
rect 74274 15940 74308 16247
rect 65649 12988 65814 13006
rect 67034 12982 67227 13265
rect 48530 7433 48720 10077
rect 44802 934 45234 7178
rect 49428 1473 49860 12133
rect 50012 7451 50180 9926
rect 53156 7403 53346 9948
rect 54054 1473 54486 12133
rect 54638 7414 54806 9969
rect 57782 7371 57972 9894
rect 58680 1473 59112 12133
rect 59264 7451 59432 10077
rect 62408 7360 62598 9926
rect 62746 7201 63178 8640
rect 63306 1473 63738 12133
rect 63890 7451 64058 9904
rect 67034 7433 67224 12982
rect 68516 12962 68687 13303
rect 69346 13354 69510 15912
rect 69346 13004 69365 13354
rect 69497 13004 69510 13354
rect 69346 12989 69510 13004
rect 70275 13356 70440 15916
rect 70275 13006 70292 13356
rect 70424 13006 70440 13356
rect 70275 12988 70440 13006
rect 71663 12982 71853 15916
rect 67372 7196 67804 10721
rect 68516 7451 68684 12962
rect 72001 12859 72433 13274
rect 73145 12962 73313 15916
rect 73971 15912 74308 15940
rect 74897 16259 75234 16286
rect 74897 15952 74926 16259
rect 75197 15952 75234 16259
rect 74897 15916 75234 15952
rect 76145 16263 76482 16286
rect 76145 15956 76177 16263
rect 76448 15956 76482 16263
rect 76145 15916 76482 15956
rect 77769 16255 78106 16286
rect 77769 15948 77800 16255
rect 78071 15948 78106 16255
rect 77769 15916 78106 15948
rect 78597 16247 78934 16282
rect 78597 15940 78629 16247
rect 78900 15940 78934 16247
rect 73972 13354 74136 15912
rect 73972 13004 73991 13354
rect 74123 13004 74136 13354
rect 73972 12989 74136 13004
rect 74901 13356 75066 15916
rect 74901 13006 74918 13356
rect 75050 13006 75066 13356
rect 74901 12988 75066 13006
rect 76289 12982 76479 15916
rect 77771 12962 77939 15916
rect 78597 15912 78934 15940
rect 79523 16259 79860 16286
rect 79523 15952 79552 16259
rect 79823 15952 79860 16259
rect 79523 15916 79860 15952
rect 80771 16263 81108 16286
rect 80771 15956 80803 16263
rect 81074 15956 81108 16263
rect 80771 15916 81108 15956
rect 82395 16255 82732 16286
rect 82395 15948 82426 16255
rect 82697 15948 82732 16255
rect 82395 15916 82732 15948
rect 83053 16247 83390 16282
rect 83053 15940 83085 16247
rect 83356 15940 83390 16247
rect 78598 13354 78762 15912
rect 78598 13004 78617 13354
rect 78749 13004 78762 13354
rect 78598 12989 78762 13004
rect 79527 13356 79692 15916
rect 79527 13006 79544 13356
rect 79676 13006 79692 13356
rect 79527 12988 79692 13006
rect 80915 12982 81105 15916
rect 82397 12962 82565 15916
rect 83053 15912 83390 15940
rect 84149 16259 84486 16286
rect 84149 15952 84178 16259
rect 84449 15952 84486 16259
rect 84149 15916 84486 15952
rect 85397 16263 85734 16286
rect 85397 15956 85429 16263
rect 85700 15956 85734 16263
rect 85397 15916 85734 15956
rect 86921 16255 87258 16286
rect 86921 15948 86952 16255
rect 87223 15948 87258 16255
rect 86921 15916 87258 15948
rect 87849 16247 88186 16282
rect 87849 15940 87881 16247
rect 88152 15940 88186 16247
rect 83224 13354 83388 15912
rect 83224 13004 83243 13354
rect 83375 13004 83388 13354
rect 83224 12989 83388 13004
rect 84153 13356 84318 15916
rect 84153 13006 84170 13356
rect 84302 13006 84318 13356
rect 84153 12988 84318 13006
rect 85541 12982 85731 15916
rect 87023 12962 87191 15916
rect 87849 15912 88186 15940
rect 88775 16259 89112 16286
rect 88775 15952 88804 16259
rect 89075 15952 89112 16259
rect 88775 15916 89112 15952
rect 90023 16263 90360 16286
rect 90023 15956 90055 16263
rect 90326 15956 90360 16263
rect 90023 15916 90360 15956
rect 91647 16255 91984 16286
rect 92505 16281 92842 16282
rect 91647 15948 91678 16255
rect 91949 15948 91984 16255
rect 91647 15916 91984 15948
rect 92476 16247 92842 16281
rect 92476 15940 92537 16247
rect 92808 15940 92842 16247
rect 87850 13354 88014 15912
rect 87850 13004 87869 13354
rect 88001 13004 88014 13354
rect 87850 12989 88014 13004
rect 88779 13356 88944 15916
rect 88779 13006 88796 13356
rect 88928 13006 88944 13356
rect 90167 13249 90357 15916
rect 91649 13287 91817 15916
rect 88779 12988 88944 13006
rect 90164 12982 90357 13249
rect 71660 7433 71850 9926
rect 67932 1461 68364 7178
rect 72558 2001 72990 12133
rect 73142 7403 73310 10023
rect 76286 7360 76476 9948
rect 77188 2001 77620 12133
rect 77768 7436 77936 10023
rect 80912 7433 81102 9937
rect 81818 2001 82250 12133
rect 82394 7446 82562 9904
rect 85538 7433 85728 9861
rect 85879 9234 86311 9811
rect 85876 7199 86308 8127
rect 86444 2001 86876 12133
rect 87020 7451 87188 9948
rect 90164 7433 90354 12982
rect 91646 12962 91817 13287
rect 92476 15912 92842 15940
rect 93401 16259 93738 16286
rect 93401 15952 93430 16259
rect 93701 15952 93738 16259
rect 93401 15916 93738 15952
rect 94649 16263 94986 16286
rect 94649 15956 94681 16263
rect 94952 15956 94986 16263
rect 94649 15916 94986 15956
rect 96073 16285 96410 16286
rect 96073 16255 96443 16285
rect 96073 15948 96104 16255
rect 96375 15948 96443 16255
rect 96073 15916 96443 15948
rect 92476 13354 92640 15912
rect 92476 13004 92495 13354
rect 92627 13004 92640 13354
rect 92476 12989 92640 13004
rect 93405 13356 93570 15916
rect 93405 13006 93422 13356
rect 93554 13006 93570 13356
rect 93405 12988 93570 13006
rect 94793 12982 94983 15916
rect 96275 12962 96443 15916
rect 97031 16247 97368 16282
rect 97031 15940 97063 16247
rect 97334 15940 97368 16247
rect 97031 15912 97368 15940
rect 98027 16259 98364 16286
rect 98027 15952 98056 16259
rect 98327 15952 98364 16259
rect 98027 15916 98364 15952
rect 98575 16263 98912 16286
rect 98575 15956 98607 16263
rect 98878 16113 98912 16263
rect 100699 16255 101036 16286
rect 101757 16281 102094 16282
rect 98878 15956 99609 16113
rect 98575 15923 99609 15956
rect 98575 15916 98912 15923
rect 97102 13354 97266 15912
rect 97102 13004 97121 13354
rect 97253 13004 97266 13354
rect 97102 12989 97266 13004
rect 98031 13356 98196 15916
rect 98031 13006 98048 13356
rect 98180 13006 98196 13356
rect 98031 12988 98196 13006
rect 99419 12982 99609 15923
rect 100699 15948 100730 16255
rect 101001 15948 101036 16255
rect 100699 15916 101036 15948
rect 101725 16247 102094 16281
rect 101725 15940 101789 16247
rect 102060 15940 102094 16247
rect 100796 15785 101069 15916
rect 100901 12962 101069 15785
rect 101725 15912 102094 15940
rect 102653 16259 102990 16286
rect 102653 15952 102682 16259
rect 102953 15952 102990 16259
rect 102653 15916 102990 15952
rect 103901 16263 104238 16286
rect 103901 15956 103933 16263
rect 104204 15956 104238 16263
rect 103901 15916 104238 15956
rect 105125 16255 105462 16286
rect 105125 15948 105156 16255
rect 105427 15948 105462 16255
rect 105125 15916 105462 15948
rect 106354 16247 106720 16282
rect 106354 15940 106415 16247
rect 106686 15940 106720 16247
rect 101725 15773 101892 15912
rect 101728 13354 101892 15773
rect 101728 13004 101747 13354
rect 101879 13004 101892 13354
rect 101728 12989 101892 13004
rect 102657 13356 102822 15916
rect 102657 13006 102674 13356
rect 102806 13006 102822 13356
rect 102657 12988 102822 13006
rect 104045 12982 104235 15916
rect 105238 15784 105695 15916
rect 105527 12962 105695 15784
rect 106354 15912 106720 15940
rect 107279 16259 107616 16286
rect 107279 15952 107308 16259
rect 107579 15952 107616 16259
rect 107279 15916 107616 15952
rect 108527 16263 108864 16286
rect 108527 15956 108559 16263
rect 108830 15956 108864 16263
rect 108527 15916 108864 15956
rect 110051 16255 110388 16286
rect 111009 16280 111346 16282
rect 110051 15948 110082 16255
rect 110353 15948 110388 16255
rect 110051 15916 110388 15948
rect 110980 16247 111346 16280
rect 110980 15940 111041 16247
rect 111312 15940 111346 16247
rect 106354 13354 106518 15912
rect 106554 15911 106718 15912
rect 106354 13004 106373 13354
rect 106505 13004 106518 13354
rect 106354 12989 106518 13004
rect 107283 13356 107448 15916
rect 107283 13006 107300 13356
rect 107432 13006 107448 13356
rect 108671 13273 108861 15916
rect 107283 12988 107448 13006
rect 108668 12982 108861 13273
rect 90502 7189 90934 10180
rect 91646 7451 91814 12962
rect 94790 7403 94980 9851
rect 95131 8730 95563 9796
rect 91070 2001 91502 7214
rect 95696 2506 96128 12019
rect 96272 7451 96440 9937
rect 99416 7433 99606 9937
rect 100322 2506 100754 11889
rect 100898 7451 101066 9850
rect 104042 7433 104232 9861
rect 104948 2506 105380 12002
rect 105524 7436 105692 9861
rect 108668 7433 108858 12982
rect 109006 7182 109438 13885
rect 110153 13287 110321 15916
rect 110150 12962 110321 13287
rect 110980 15912 111346 15940
rect 111905 16259 112242 16286
rect 111905 15952 111934 16259
rect 112205 15952 112242 16259
rect 111905 15916 112242 15952
rect 113153 16263 113490 16286
rect 113153 15956 113185 16263
rect 113456 15956 113490 16263
rect 113153 15916 113490 15956
rect 114777 16255 115114 16286
rect 114777 15948 114808 16255
rect 115079 15948 115114 16255
rect 114777 15916 115114 15948
rect 115606 16247 115972 16282
rect 115606 15940 115667 16247
rect 115938 15940 115972 16247
rect 110980 13354 111144 15912
rect 110980 13004 110999 13354
rect 111131 13004 111144 13354
rect 110980 12989 111144 13004
rect 111909 13356 112074 15916
rect 111909 13006 111926 13356
rect 112058 13006 112074 13356
rect 111909 12988 112074 13006
rect 113297 12982 113487 15916
rect 114779 12962 114947 15916
rect 115606 15912 115972 15940
rect 116531 16259 116868 16286
rect 116531 15952 116560 16259
rect 116831 15952 116868 16259
rect 116531 15916 116868 15952
rect 117779 16263 118116 16286
rect 117779 15956 117811 16263
rect 118082 15956 118116 16263
rect 117779 15916 118116 15956
rect 119303 16255 119640 16286
rect 119303 15948 119334 16255
rect 119605 15948 119640 16255
rect 119303 15916 119640 15948
rect 120232 16282 120396 16287
rect 120232 16247 120598 16282
rect 120232 15940 120293 16247
rect 120564 15940 120598 16247
rect 115606 13354 115770 15912
rect 115606 13004 115625 13354
rect 115757 13004 115770 13354
rect 115606 12989 115770 13004
rect 116535 13356 116700 15916
rect 116535 13006 116552 13356
rect 116684 13006 116700 13356
rect 116535 12988 116700 13006
rect 117923 12982 118113 15916
rect 119405 12962 119573 15916
rect 120232 15912 120598 15940
rect 121157 16259 121494 16286
rect 121157 15952 121186 16259
rect 121457 15952 121494 16259
rect 121157 15916 121494 15952
rect 122405 16263 122742 16286
rect 122405 15956 122437 16263
rect 122708 15956 122742 16263
rect 122405 15916 122742 15956
rect 124029 16255 124366 16286
rect 124029 15948 124060 16255
rect 124331 15948 124366 16255
rect 124029 15916 124366 15948
rect 124858 16282 125033 16283
rect 124858 16247 125224 16282
rect 124858 15940 124919 16247
rect 125190 15940 125224 16247
rect 120232 13354 120396 15912
rect 120232 13004 120251 13354
rect 120383 13004 120396 13354
rect 120232 12989 120396 13004
rect 121161 13356 121326 15916
rect 121161 13006 121178 13356
rect 121310 13006 121326 13356
rect 122549 13265 122739 15916
rect 124031 13303 124199 15916
rect 121161 12988 121326 13006
rect 122546 12982 122739 13265
rect 110150 7451 110318 12962
rect 113294 7433 113484 9948
rect 113635 9239 114067 9811
rect 109574 2506 110006 7226
rect 114200 4617 114632 11997
rect 114776 7436 114944 9904
rect 117920 7433 118110 9883
rect 118826 4617 119258 11996
rect 119402 7414 119570 9883
rect 122546 7433 122736 12982
rect 124028 12962 124199 13303
rect 124858 15912 125224 15940
rect 125783 16259 126120 16286
rect 125783 15952 125812 16259
rect 126083 15952 126120 16259
rect 125783 15916 126120 15952
rect 127031 16263 127368 16286
rect 127031 15956 127063 16263
rect 127334 15956 127368 16263
rect 127031 15916 127368 15956
rect 128455 16285 128792 16286
rect 128455 16255 128825 16285
rect 128455 15948 128486 16255
rect 128757 15948 128825 16255
rect 128455 15916 128825 15948
rect 124858 15737 125033 15912
rect 124858 13354 125022 15737
rect 124858 13004 124877 13354
rect 125009 13004 125022 13354
rect 124858 12989 125022 13004
rect 125787 13356 125952 15916
rect 125787 13006 125804 13356
rect 125936 13006 125952 13356
rect 125787 12988 125952 13006
rect 127175 12982 127365 15916
rect 128657 12962 128825 15916
rect 129484 16282 129648 16283
rect 129484 16247 129850 16282
rect 129484 15940 129545 16247
rect 129816 15940 129850 16247
rect 129484 15912 129850 15940
rect 130409 16259 130746 16286
rect 130409 15952 130438 16259
rect 130709 15952 130746 16259
rect 130409 15916 130746 15952
rect 131657 16263 131994 16286
rect 131657 15956 131689 16263
rect 131960 15956 131994 16263
rect 131657 15916 131994 15956
rect 133281 16255 133618 16286
rect 134110 16282 134274 16283
rect 133281 15948 133312 16255
rect 133583 15948 133618 16255
rect 133281 15916 133618 15948
rect 133839 16247 134274 16282
rect 133839 15940 133871 16247
rect 134142 15940 134274 16247
rect 129484 13354 129648 15912
rect 129484 13004 129503 13354
rect 129635 13004 129648 13354
rect 129484 12989 129648 13004
rect 130413 13356 130578 15916
rect 130413 13006 130430 13356
rect 130562 13006 130578 13356
rect 130413 12988 130578 13006
rect 131801 12982 131991 15916
rect 133283 12962 133451 15916
rect 133839 15912 134274 15940
rect 135035 16259 135372 16286
rect 135035 15952 135064 16259
rect 135335 15952 135372 16259
rect 135035 15916 135372 15952
rect 136283 16263 136620 16286
rect 136283 15956 136315 16263
rect 136586 15956 136620 16263
rect 136283 15916 136620 15956
rect 137907 16255 138244 16286
rect 137907 15948 137938 16255
rect 138209 15948 138244 16255
rect 137907 15916 138244 15948
rect 134110 13314 134274 15912
rect 134110 12964 134129 13314
rect 134261 12964 134274 13314
rect 124028 7451 124196 12962
rect 134110 12949 134274 12964
rect 135039 13316 135204 15916
rect 135039 12966 135056 13316
rect 135188 12966 135204 13316
rect 136427 13273 136617 15916
rect 137909 13287 138077 15916
rect 135039 12948 135204 12966
rect 136424 12982 136617 13273
rect 127172 7414 127362 9937
rect 128078 4617 128510 12052
rect 128654 7403 128822 9980
rect 131798 7433 131988 9840
rect 132704 4617 133136 12037
rect 133280 7349 133448 9883
rect 136424 7433 136614 12982
rect 137906 12962 138077 13287
rect 137326 7203 137758 7638
rect 137906 7451 138074 12962
<< via2 >>
rect -183 15940 88 16247
rect 910 15952 1181 16259
rect 2161 15956 2432 16263
rect 3784 15948 4055 16255
rect 4443 15940 4714 16247
rect 5536 15952 5807 16259
rect 6787 15956 7058 16263
rect 8410 15948 8681 16255
rect 9069 15940 9340 16247
rect 10162 15952 10433 16259
rect 11413 15956 11684 16263
rect 13036 15948 13307 16255
rect 13895 15940 14166 16247
rect 14788 15952 15059 16259
rect 16039 15956 16310 16263
rect 17662 15948 17933 16255
rect 18321 15940 18592 16247
rect 19414 15952 19685 16259
rect 20665 15956 20936 16263
rect 22288 15948 22559 16255
rect 22947 15940 23218 16247
rect 24040 15952 24311 16259
rect 25601 15956 25872 16263
rect 26314 15948 26585 16255
rect 27513 15940 27784 16247
rect 28766 15952 29037 16259
rect 29917 15956 30188 16263
rect 31540 15948 31811 16255
rect 32199 15940 32470 16247
rect 33292 15952 33563 16259
rect 34543 15956 34814 16263
rect 36166 15948 36437 16255
rect 36825 15940 37096 16247
rect 37918 15952 38189 16259
rect 39169 15956 39440 16263
rect 40792 15948 41063 16255
rect 41451 15940 41722 16247
rect 42544 15952 42815 16259
rect 43795 15956 44066 16263
rect 45418 15948 45689 16255
rect 46077 15940 46348 16247
rect 47170 15952 47441 16259
rect 48421 15956 48692 16263
rect 50044 15948 50315 16255
rect 50703 15940 50974 16247
rect 51796 15952 52067 16259
rect 53047 15956 53318 16263
rect 54670 15948 54941 16255
rect 55329 15940 55600 16247
rect 56422 15952 56693 16259
rect 57673 15956 57944 16263
rect 59296 15948 59567 16255
rect 59955 15940 60226 16247
rect 61048 15952 61319 16259
rect 61899 15956 62170 16263
rect 64222 15948 64493 16255
rect 64881 15940 65152 16247
rect 65674 15952 65945 16259
rect 67106 15956 67377 16263
rect 68548 15948 68819 16255
rect 69207 15940 69478 16247
rect 70300 15952 70571 16259
rect 71551 15956 71822 16263
rect 73174 15948 73445 16255
rect 74003 15940 74274 16247
rect 74926 15952 75197 16259
rect 76177 15956 76448 16263
rect 77800 15948 78071 16255
rect 78629 15940 78900 16247
rect 79552 15952 79823 16259
rect 80803 15956 81074 16263
rect 82426 15948 82697 16255
rect 83085 15940 83356 16247
rect 84178 15952 84449 16259
rect 85429 15956 85700 16263
rect 86952 15948 87223 16255
rect 87881 15940 88152 16247
rect 88804 15952 89075 16259
rect 90055 15956 90326 16263
rect 91678 15948 91949 16255
rect 92537 15940 92808 16247
rect 93430 15952 93701 16259
rect 94681 15956 94952 16263
rect 96104 15948 96375 16255
rect 97063 15940 97334 16247
rect 98056 15952 98327 16259
rect 98607 15956 98878 16263
rect 100730 15948 101001 16255
rect 101789 15940 102060 16247
rect 102682 15952 102953 16259
rect 103933 15956 104204 16263
rect 105156 15948 105427 16255
rect 106415 15940 106686 16247
rect 107308 15952 107579 16259
rect 108559 15956 108830 16263
rect 110082 15948 110353 16255
rect 111041 15940 111312 16247
rect 111934 15952 112205 16259
rect 113185 15956 113456 16263
rect 114808 15948 115079 16255
rect 115667 15940 115938 16247
rect 116560 15952 116831 16259
rect 117811 15956 118082 16263
rect 119334 15948 119605 16255
rect 120293 15940 120564 16247
rect 121186 15952 121457 16259
rect 122437 15956 122708 16263
rect 124060 15948 124331 16255
rect 124919 15940 125190 16247
rect 125812 15952 126083 16259
rect 127063 15956 127334 16263
rect 128486 15948 128757 16255
rect 129545 15940 129816 16247
rect 130438 15952 130709 16259
rect 131689 15956 131960 16263
rect 133312 15948 133583 16255
rect 133871 15940 134142 16247
rect 135064 15952 135335 16259
rect 136315 15956 136586 16263
rect 137938 15948 138209 16255
<< metal3 >>
rect -215 16247 122 16282
rect -215 15940 -183 16247
rect 88 15940 122 16247
rect -215 15912 122 15940
rect 881 16259 1218 16286
rect 881 15952 910 16259
rect 1181 15952 1218 16259
rect 881 15916 1218 15952
rect 2129 16263 2466 16286
rect 2129 15956 2161 16263
rect 2432 15956 2466 16263
rect 2129 15916 2466 15956
rect 3753 16255 4090 16286
rect 3753 15948 3784 16255
rect 4055 15948 4090 16255
rect 3753 15916 4090 15948
rect 4411 16247 4748 16282
rect 4411 15940 4443 16247
rect 4714 15940 4748 16247
rect 4411 15912 4748 15940
rect 5507 16259 5844 16286
rect 5507 15952 5536 16259
rect 5807 15952 5844 16259
rect 5507 15916 5844 15952
rect 6755 16263 7092 16286
rect 6755 15956 6787 16263
rect 7058 15956 7092 16263
rect 6755 15916 7092 15956
rect 8379 16255 8716 16286
rect 8379 15948 8410 16255
rect 8681 15948 8716 16255
rect 8379 15916 8716 15948
rect 9037 16247 9374 16282
rect 9037 15940 9069 16247
rect 9340 15940 9374 16247
rect 9037 15912 9374 15940
rect 10133 16259 10470 16286
rect 10133 15952 10162 16259
rect 10433 15952 10470 16259
rect 10133 15916 10470 15952
rect 11381 16263 11718 16286
rect 11381 15956 11413 16263
rect 11684 15956 11718 16263
rect 11381 15916 11718 15956
rect 13005 16255 13342 16286
rect 13005 15948 13036 16255
rect 13307 15948 13342 16255
rect 13005 15916 13342 15948
rect 13863 16247 14200 16282
rect 13863 15940 13895 16247
rect 14166 15940 14200 16247
rect 13863 15912 14200 15940
rect 14759 16259 15096 16286
rect 14759 15952 14788 16259
rect 15059 15952 15096 16259
rect 14759 15916 15096 15952
rect 16007 16263 16344 16286
rect 16007 15956 16039 16263
rect 16310 15956 16344 16263
rect 16007 15916 16344 15956
rect 17631 16255 17968 16286
rect 17631 15948 17662 16255
rect 17933 15948 17968 16255
rect 17631 15916 17968 15948
rect 18289 16247 18626 16282
rect 18289 15940 18321 16247
rect 18592 15940 18626 16247
rect 18289 15912 18626 15940
rect 19385 16259 19722 16286
rect 19385 15952 19414 16259
rect 19685 15952 19722 16259
rect 19385 15916 19722 15952
rect 20633 16263 20970 16286
rect 20633 15956 20665 16263
rect 20936 15956 20970 16263
rect 20633 15916 20970 15956
rect 22257 16255 22594 16286
rect 22257 15948 22288 16255
rect 22559 15948 22594 16255
rect 22257 15916 22594 15948
rect 22915 16247 23252 16282
rect 22915 15940 22947 16247
rect 23218 15940 23252 16247
rect 22915 15912 23252 15940
rect 24011 16259 24348 16286
rect 24011 15952 24040 16259
rect 24311 15952 24348 16259
rect 24011 15916 24348 15952
rect 25569 16263 25906 16286
rect 25569 15956 25601 16263
rect 25872 15956 25906 16263
rect 25569 15916 25906 15956
rect 26283 16255 26620 16286
rect 26283 15948 26314 16255
rect 26585 15948 26620 16255
rect 26283 15916 26620 15948
rect 27481 16247 27818 16282
rect 27481 15940 27513 16247
rect 27784 15940 27818 16247
rect 27481 15912 27818 15940
rect 28737 16259 29074 16286
rect 28737 15952 28766 16259
rect 29037 15952 29074 16259
rect 28737 15916 29074 15952
rect 29885 16263 30222 16286
rect 29885 15956 29917 16263
rect 30188 15956 30222 16263
rect 29885 15916 30222 15956
rect 31509 16255 31846 16286
rect 31509 15948 31540 16255
rect 31811 15948 31846 16255
rect 31509 15916 31846 15948
rect 32167 16247 32504 16282
rect 32167 15940 32199 16247
rect 32470 15940 32504 16247
rect 32167 15912 32504 15940
rect 33263 16259 33600 16286
rect 33263 15952 33292 16259
rect 33563 15952 33600 16259
rect 33263 15916 33600 15952
rect 34511 16263 34848 16286
rect 34511 15956 34543 16263
rect 34814 15956 34848 16263
rect 34511 15916 34848 15956
rect 36135 16255 36472 16286
rect 36135 15948 36166 16255
rect 36437 15948 36472 16255
rect 36135 15916 36472 15948
rect 36793 16247 37130 16282
rect 36793 15940 36825 16247
rect 37096 15940 37130 16247
rect 36793 15912 37130 15940
rect 37889 16259 38226 16286
rect 37889 15952 37918 16259
rect 38189 15952 38226 16259
rect 37889 15916 38226 15952
rect 39137 16263 39474 16286
rect 39137 15956 39169 16263
rect 39440 15956 39474 16263
rect 39137 15916 39474 15956
rect 40761 16255 41098 16286
rect 40761 15948 40792 16255
rect 41063 15948 41098 16255
rect 40761 15916 41098 15948
rect 41419 16247 41756 16282
rect 41419 15940 41451 16247
rect 41722 15940 41756 16247
rect 41419 15912 41756 15940
rect 42515 16259 42852 16286
rect 42515 15952 42544 16259
rect 42815 15952 42852 16259
rect 42515 15916 42852 15952
rect 43763 16263 44100 16286
rect 43763 15956 43795 16263
rect 44066 15956 44100 16263
rect 43763 15916 44100 15956
rect 45387 16255 45724 16286
rect 45387 15948 45418 16255
rect 45689 15948 45724 16255
rect 45387 15916 45724 15948
rect 46045 16247 46382 16282
rect 46045 15940 46077 16247
rect 46348 15940 46382 16247
rect 46045 15912 46382 15940
rect 47141 16259 47478 16286
rect 47141 15952 47170 16259
rect 47441 15952 47478 16259
rect 47141 15916 47478 15952
rect 48389 16263 48726 16286
rect 48389 15956 48421 16263
rect 48692 15956 48726 16263
rect 48389 15916 48726 15956
rect 50013 16255 50350 16286
rect 50013 15948 50044 16255
rect 50315 15948 50350 16255
rect 50013 15916 50350 15948
rect 50671 16247 51008 16282
rect 50671 15940 50703 16247
rect 50974 15940 51008 16247
rect 50671 15912 51008 15940
rect 51767 16259 52104 16286
rect 51767 15952 51796 16259
rect 52067 15952 52104 16259
rect 51767 15916 52104 15952
rect 53015 16263 53352 16286
rect 53015 15956 53047 16263
rect 53318 15956 53352 16263
rect 53015 15916 53352 15956
rect 54639 16255 54976 16286
rect 54639 15948 54670 16255
rect 54941 15948 54976 16255
rect 54639 15916 54976 15948
rect 55297 16247 55634 16282
rect 55297 15940 55329 16247
rect 55600 15940 55634 16247
rect 55297 15912 55634 15940
rect 56393 16259 56730 16286
rect 56393 15952 56422 16259
rect 56693 15952 56730 16259
rect 56393 15916 56730 15952
rect 57641 16263 57978 16286
rect 57641 15956 57673 16263
rect 57944 15956 57978 16263
rect 57641 15916 57978 15956
rect 59265 16255 59602 16286
rect 59265 15948 59296 16255
rect 59567 15948 59602 16255
rect 59265 15916 59602 15948
rect 59923 16247 60260 16282
rect 59923 15940 59955 16247
rect 60226 15940 60260 16247
rect 59923 15912 60260 15940
rect 61019 16259 61356 16286
rect 61019 15952 61048 16259
rect 61319 15952 61356 16259
rect 61019 15916 61356 15952
rect 61867 16263 62204 16286
rect 61867 15956 61899 16263
rect 62170 15956 62204 16263
rect 61867 15916 62204 15956
rect 64191 16255 64528 16286
rect 64191 15948 64222 16255
rect 64493 15948 64528 16255
rect 64191 15916 64528 15948
rect 64849 16247 65186 16282
rect 64849 15940 64881 16247
rect 65152 15940 65186 16247
rect 64849 15912 65186 15940
rect 65645 16259 65982 16286
rect 65645 15952 65674 16259
rect 65945 15952 65982 16259
rect 65645 15916 65982 15952
rect 67074 16263 67411 16286
rect 67074 15956 67106 16263
rect 67377 15956 67411 16263
rect 67074 15916 67411 15956
rect 68517 16255 68854 16286
rect 68517 15948 68548 16255
rect 68819 15948 68854 16255
rect 68517 15916 68854 15948
rect 69175 16247 69512 16282
rect 69175 15940 69207 16247
rect 69478 15940 69512 16247
rect 69175 15912 69512 15940
rect 70271 16259 70608 16286
rect 70271 15952 70300 16259
rect 70571 15952 70608 16259
rect 70271 15916 70608 15952
rect 71519 16263 71856 16286
rect 71519 15956 71551 16263
rect 71822 15956 71856 16263
rect 71519 15916 71856 15956
rect 73143 16255 73480 16286
rect 73143 15948 73174 16255
rect 73445 15948 73480 16255
rect 73143 15916 73480 15948
rect 73971 16247 74308 16282
rect 73971 15940 74003 16247
rect 74274 15940 74308 16247
rect 73971 15912 74308 15940
rect 74897 16259 75234 16286
rect 74897 15952 74926 16259
rect 75197 15952 75234 16259
rect 74897 15916 75234 15952
rect 76145 16263 76482 16286
rect 76145 15956 76177 16263
rect 76448 15956 76482 16263
rect 76145 15916 76482 15956
rect 77769 16255 78106 16286
rect 77769 15948 77800 16255
rect 78071 15948 78106 16255
rect 77769 15916 78106 15948
rect 78597 16247 78934 16282
rect 78597 15940 78629 16247
rect 78900 15940 78934 16247
rect 78597 15912 78934 15940
rect 79523 16259 79860 16286
rect 79523 15952 79552 16259
rect 79823 15952 79860 16259
rect 79523 15916 79860 15952
rect 80771 16263 81108 16286
rect 80771 15956 80803 16263
rect 81074 15956 81108 16263
rect 80771 15916 81108 15956
rect 82395 16255 82732 16286
rect 82395 15948 82426 16255
rect 82697 15948 82732 16255
rect 82395 15916 82732 15948
rect 83053 16247 83390 16282
rect 83053 15940 83085 16247
rect 83356 15940 83390 16247
rect 83053 15912 83390 15940
rect 84149 16259 84486 16286
rect 84149 15952 84178 16259
rect 84449 15952 84486 16259
rect 84149 15916 84486 15952
rect 85397 16263 85734 16286
rect 85397 15956 85429 16263
rect 85700 15956 85734 16263
rect 85397 15916 85734 15956
rect 86921 16255 87258 16286
rect 86921 15948 86952 16255
rect 87223 15948 87258 16255
rect 86921 15916 87258 15948
rect 87849 16247 88186 16282
rect 87849 15940 87881 16247
rect 88152 15940 88186 16247
rect 87849 15912 88186 15940
rect 88775 16259 89112 16286
rect 88775 15952 88804 16259
rect 89075 15952 89112 16259
rect 88775 15916 89112 15952
rect 90023 16263 90360 16286
rect 90023 15956 90055 16263
rect 90326 15956 90360 16263
rect 90023 15916 90360 15956
rect 91647 16255 91984 16286
rect 91647 15948 91678 16255
rect 91949 15948 91984 16255
rect 91647 15916 91984 15948
rect 92505 16247 92842 16282
rect 92505 15940 92537 16247
rect 92808 15940 92842 16247
rect 92505 15912 92842 15940
rect 93401 16259 93738 16286
rect 93401 15952 93430 16259
rect 93701 15952 93738 16259
rect 93401 15916 93738 15952
rect 94649 16263 94986 16286
rect 94649 15956 94681 16263
rect 94952 15956 94986 16263
rect 94649 15916 94986 15956
rect 96073 16255 96410 16286
rect 96073 15948 96104 16255
rect 96375 15948 96410 16255
rect 96073 15916 96410 15948
rect 97031 16247 97368 16282
rect 97031 15940 97063 16247
rect 97334 15940 97368 16247
rect 97031 15912 97368 15940
rect 98027 16259 98364 16286
rect 98027 15952 98056 16259
rect 98327 15952 98364 16259
rect 98027 15916 98364 15952
rect 98575 16263 98912 16286
rect 98575 15956 98607 16263
rect 98878 15956 98912 16263
rect 98575 15916 98912 15956
rect 100699 16255 101036 16286
rect 100699 15948 100730 16255
rect 101001 15948 101036 16255
rect 100699 15916 101036 15948
rect 101757 16247 102094 16282
rect 101757 15940 101789 16247
rect 102060 15940 102094 16247
rect 101757 15912 102094 15940
rect 102653 16259 102990 16286
rect 102653 15952 102682 16259
rect 102953 15952 102990 16259
rect 102653 15916 102990 15952
rect 103901 16263 104238 16286
rect 103901 15956 103933 16263
rect 104204 15956 104238 16263
rect 103901 15916 104238 15956
rect 105125 16255 105462 16286
rect 105125 15948 105156 16255
rect 105427 15948 105462 16255
rect 105125 15916 105462 15948
rect 106383 16247 106720 16282
rect 106383 15940 106415 16247
rect 106686 15940 106720 16247
rect 106383 15912 106720 15940
rect 107279 16259 107616 16286
rect 107279 15952 107308 16259
rect 107579 15952 107616 16259
rect 107279 15916 107616 15952
rect 108527 16263 108864 16286
rect 108527 15956 108559 16263
rect 108830 15956 108864 16263
rect 108527 15916 108864 15956
rect 110051 16255 110388 16286
rect 110051 15948 110082 16255
rect 110353 15948 110388 16255
rect 110051 15916 110388 15948
rect 111009 16247 111346 16282
rect 111009 15940 111041 16247
rect 111312 15940 111346 16247
rect 111009 15912 111346 15940
rect 111905 16259 112242 16286
rect 111905 15952 111934 16259
rect 112205 15952 112242 16259
rect 111905 15916 112242 15952
rect 113153 16263 113490 16286
rect 113153 15956 113185 16263
rect 113456 15956 113490 16263
rect 113153 15916 113490 15956
rect 114777 16255 115114 16286
rect 114777 15948 114808 16255
rect 115079 15948 115114 16255
rect 114777 15916 115114 15948
rect 115635 16247 115972 16282
rect 115635 15940 115667 16247
rect 115938 15940 115972 16247
rect 115635 15912 115972 15940
rect 116531 16259 116868 16286
rect 116531 15952 116560 16259
rect 116831 15952 116868 16259
rect 116531 15916 116868 15952
rect 117779 16263 118116 16286
rect 117779 15956 117811 16263
rect 118082 15956 118116 16263
rect 117779 15916 118116 15956
rect 119303 16255 119640 16286
rect 119303 15948 119334 16255
rect 119605 15948 119640 16255
rect 119303 15916 119640 15948
rect 120261 16247 120598 16282
rect 120261 15940 120293 16247
rect 120564 15940 120598 16247
rect 120261 15912 120598 15940
rect 121157 16259 121494 16286
rect 121157 15952 121186 16259
rect 121457 15952 121494 16259
rect 121157 15916 121494 15952
rect 122405 16263 122742 16286
rect 122405 15956 122437 16263
rect 122708 15956 122742 16263
rect 122405 15916 122742 15956
rect 124029 16255 124366 16286
rect 124029 15948 124060 16255
rect 124331 15948 124366 16255
rect 124029 15916 124366 15948
rect 124887 16247 125224 16282
rect 124887 15940 124919 16247
rect 125190 15940 125224 16247
rect 124887 15912 125224 15940
rect 125783 16259 126120 16286
rect 125783 15952 125812 16259
rect 126083 15952 126120 16259
rect 125783 15916 126120 15952
rect 127031 16263 127368 16286
rect 127031 15956 127063 16263
rect 127334 15956 127368 16263
rect 127031 15916 127368 15956
rect 128455 16255 128792 16286
rect 128455 15948 128486 16255
rect 128757 15948 128792 16255
rect 128455 15916 128792 15948
rect 129513 16247 129850 16282
rect 129513 15940 129545 16247
rect 129816 15940 129850 16247
rect 129513 15912 129850 15940
rect 130409 16259 130746 16286
rect 130409 15952 130438 16259
rect 130709 15952 130746 16259
rect 130409 15916 130746 15952
rect 131657 16263 131994 16286
rect 131657 15956 131689 16263
rect 131960 15956 131994 16263
rect 131657 15916 131994 15956
rect 133281 16255 133618 16286
rect 133281 15948 133312 16255
rect 133583 15948 133618 16255
rect 133281 15916 133618 15948
rect 133839 16247 134176 16282
rect 133839 15940 133871 16247
rect 134142 15940 134176 16247
rect 133839 15912 134176 15940
rect 135035 16259 135372 16286
rect 135035 15952 135064 16259
rect 135335 15952 135372 16259
rect 135035 15916 135372 15952
rect 136283 16263 136620 16286
rect 136283 15956 136315 16263
rect 136586 15956 136620 16263
rect 136283 15916 136620 15956
rect 137907 16255 138244 16286
rect 137907 15948 137938 16255
rect 138209 15948 138244 16255
rect 137907 15916 138244 15948
rect -80 13751 140525 13879
rect -80 13239 140525 13367
rect -80 12727 140525 12855
rect -80 12215 140525 12343
rect -80 11703 140525 11831
rect -80 11191 140525 11319
rect -80 10679 140525 10807
rect -80 10167 140525 10295
rect -80 9655 140525 9783
rect -80 9143 140525 9271
rect -80 8631 140525 8759
rect -80 8119 140525 8247
rect -80 7607 140525 7735
rect -80 7095 140525 7223
rect -80 6583 140525 6711
rect -80 6071 140525 6199
rect -80 5559 140525 5687
rect -80 5047 140525 5175
rect -80 4535 140525 4663
rect -80 4023 140525 4151
rect -80 2487 140525 2615
rect -80 1975 140525 2103
rect -80 1463 140525 1591
rect -80 951 140525 1079
rect -80 439 140525 567
<< via3 >>
rect -183 15940 88 16247
rect 910 15952 1181 16259
rect 2161 15956 2432 16263
rect 3784 15948 4055 16255
rect 4443 15940 4714 16247
rect 5536 15952 5807 16259
rect 6787 15956 7058 16263
rect 8410 15948 8681 16255
rect 9069 15940 9340 16247
rect 10162 15952 10433 16259
rect 11413 15956 11684 16263
rect 13036 15948 13307 16255
rect 13895 15940 14166 16247
rect 14788 15952 15059 16259
rect 16039 15956 16310 16263
rect 17662 15948 17933 16255
rect 18321 15940 18592 16247
rect 19414 15952 19685 16259
rect 20665 15956 20936 16263
rect 22288 15948 22559 16255
rect 22947 15940 23218 16247
rect 24040 15952 24311 16259
rect 25601 15956 25872 16263
rect 26314 15948 26585 16255
rect 27513 15940 27784 16247
rect 28766 15952 29037 16259
rect 29917 15956 30188 16263
rect 31540 15948 31811 16255
rect 32199 15940 32470 16247
rect 33292 15952 33563 16259
rect 34543 15956 34814 16263
rect 36166 15948 36437 16255
rect 36825 15940 37096 16247
rect 37918 15952 38189 16259
rect 39169 15956 39440 16263
rect 40792 15948 41063 16255
rect 41451 15940 41722 16247
rect 42544 15952 42815 16259
rect 43795 15956 44066 16263
rect 45418 15948 45689 16255
rect 46077 15940 46348 16247
rect 47170 15952 47441 16259
rect 48421 15956 48692 16263
rect 50044 15948 50315 16255
rect 50703 15940 50974 16247
rect 51796 15952 52067 16259
rect 53047 15956 53318 16263
rect 54670 15948 54941 16255
rect 55329 15940 55600 16247
rect 56422 15952 56693 16259
rect 57673 15956 57944 16263
rect 59296 15948 59567 16255
rect 59955 15940 60226 16247
rect 61048 15952 61319 16259
rect 61899 15956 62170 16263
rect 64222 15948 64493 16255
rect 64881 15940 65152 16247
rect 65674 15952 65945 16259
rect 67106 15956 67377 16263
rect 68548 15948 68819 16255
rect 69207 15940 69478 16247
rect 70300 15952 70571 16259
rect 71551 15956 71822 16263
rect 73174 15948 73445 16255
rect 74003 15940 74274 16247
rect 74926 15952 75197 16259
rect 76177 15956 76448 16263
rect 77800 15948 78071 16255
rect 78629 15940 78900 16247
rect 79552 15952 79823 16259
rect 80803 15956 81074 16263
rect 82426 15948 82697 16255
rect 83085 15940 83356 16247
rect 84178 15952 84449 16259
rect 85429 15956 85700 16263
rect 86952 15948 87223 16255
rect 87881 15940 88152 16247
rect 88804 15952 89075 16259
rect 90055 15956 90326 16263
rect 91678 15948 91949 16255
rect 92537 15940 92808 16247
rect 93430 15952 93701 16259
rect 94681 15956 94952 16263
rect 96104 15948 96375 16255
rect 97063 15940 97334 16247
rect 98056 15952 98327 16259
rect 98607 15956 98878 16263
rect 100730 15948 101001 16255
rect 101789 15940 102060 16247
rect 102682 15952 102953 16259
rect 103933 15956 104204 16263
rect 105156 15948 105427 16255
rect 106415 15940 106686 16247
rect 107308 15952 107579 16259
rect 108559 15956 108830 16263
rect 110082 15948 110353 16255
rect 111041 15940 111312 16247
rect 111934 15952 112205 16259
rect 113185 15956 113456 16263
rect 114808 15948 115079 16255
rect 115667 15940 115938 16247
rect 116560 15952 116831 16259
rect 117811 15956 118082 16263
rect 119334 15948 119605 16255
rect 120293 15940 120564 16247
rect 121186 15952 121457 16259
rect 122437 15956 122708 16263
rect 124060 15948 124331 16255
rect 124919 15940 125190 16247
rect 125812 15952 126083 16259
rect 127063 15956 127334 16263
rect 128486 15948 128757 16255
rect 129545 15940 129816 16247
rect 130438 15952 130709 16259
rect 131689 15956 131960 16263
rect 133312 15948 133583 16255
rect 133871 15940 134142 16247
rect 135064 15952 135335 16259
rect 136315 15956 136586 16263
rect 137938 15948 138209 16255
<< metal4 >>
rect -215 16247 122 16282
rect -215 15940 -183 16247
rect 88 15940 122 16247
rect -215 15912 122 15940
rect 881 16259 1218 16286
rect 881 15952 910 16259
rect 1181 15952 1218 16259
rect 881 15916 1218 15952
rect 2129 16263 2466 16286
rect 2129 15956 2161 16263
rect 2432 15956 2466 16263
rect 2129 15916 2466 15956
rect 3753 16255 4090 16286
rect 3753 15948 3784 16255
rect 4055 15948 4090 16255
rect 3753 15916 4090 15948
rect 4411 16247 4748 16282
rect 4411 15940 4443 16247
rect 4714 15940 4748 16247
rect 4411 15912 4748 15940
rect 5507 16259 5844 16286
rect 5507 15952 5536 16259
rect 5807 15952 5844 16259
rect 5507 15916 5844 15952
rect 6755 16263 7092 16286
rect 6755 15956 6787 16263
rect 7058 15956 7092 16263
rect 6755 15916 7092 15956
rect 8379 16255 8716 16286
rect 8379 15948 8410 16255
rect 8681 15948 8716 16255
rect 8379 15916 8716 15948
rect 9037 16247 9374 16282
rect 9037 15940 9069 16247
rect 9340 15940 9374 16247
rect 9037 15912 9374 15940
rect 10133 16259 10470 16286
rect 10133 15952 10162 16259
rect 10433 15952 10470 16259
rect 10133 15916 10470 15952
rect 11381 16263 11718 16286
rect 11381 15956 11413 16263
rect 11684 15956 11718 16263
rect 11381 15916 11718 15956
rect 13005 16255 13342 16286
rect 13005 15948 13036 16255
rect 13307 15948 13342 16255
rect 13005 15916 13342 15948
rect 13863 16247 14200 16282
rect 13863 15940 13895 16247
rect 14166 15940 14200 16247
rect 13863 15912 14200 15940
rect 14759 16259 15096 16286
rect 14759 15952 14788 16259
rect 15059 15952 15096 16259
rect 14759 15916 15096 15952
rect 16007 16263 16344 16286
rect 16007 15956 16039 16263
rect 16310 15956 16344 16263
rect 16007 15916 16344 15956
rect 17631 16255 17968 16286
rect 17631 15948 17662 16255
rect 17933 15948 17968 16255
rect 17631 15916 17968 15948
rect 18289 16247 18626 16282
rect 18289 15940 18321 16247
rect 18592 15940 18626 16247
rect 18289 15912 18626 15940
rect 19385 16259 19722 16286
rect 19385 15952 19414 16259
rect 19685 15952 19722 16259
rect 19385 15916 19722 15952
rect 20633 16263 20970 16286
rect 20633 15956 20665 16263
rect 20936 15956 20970 16263
rect 20633 15916 20970 15956
rect 22257 16255 22594 16286
rect 22257 15948 22288 16255
rect 22559 15948 22594 16255
rect 22257 15916 22594 15948
rect 22915 16247 23252 16282
rect 22915 15940 22947 16247
rect 23218 15940 23252 16247
rect 22915 15912 23252 15940
rect 24011 16259 24348 16286
rect 24011 15952 24040 16259
rect 24311 15952 24348 16259
rect 24011 15916 24348 15952
rect 25569 16263 25906 16286
rect 25569 15956 25601 16263
rect 25872 15956 25906 16263
rect 25569 15916 25906 15956
rect 26283 16255 26620 16286
rect 26283 15948 26314 16255
rect 26585 15948 26620 16255
rect 26283 15916 26620 15948
rect 27481 16247 27818 16282
rect 27481 15940 27513 16247
rect 27784 15940 27818 16247
rect 27481 15912 27818 15940
rect 28737 16259 29074 16286
rect 28737 15952 28766 16259
rect 29037 15952 29074 16259
rect 28737 15916 29074 15952
rect 29885 16263 30222 16286
rect 29885 15956 29917 16263
rect 30188 15956 30222 16263
rect 29885 15916 30222 15956
rect 31509 16255 31846 16286
rect 31509 15948 31540 16255
rect 31811 15948 31846 16255
rect 31509 15916 31846 15948
rect 32167 16247 32504 16282
rect 32167 15940 32199 16247
rect 32470 15940 32504 16247
rect 32167 15912 32504 15940
rect 33263 16259 33600 16286
rect 33263 15952 33292 16259
rect 33563 15952 33600 16259
rect 33263 15916 33600 15952
rect 34511 16263 34848 16286
rect 34511 15956 34543 16263
rect 34814 15956 34848 16263
rect 34511 15916 34848 15956
rect 36135 16255 36472 16286
rect 36135 15948 36166 16255
rect 36437 15948 36472 16255
rect 36135 15916 36472 15948
rect 36793 16247 37130 16282
rect 36793 15940 36825 16247
rect 37096 15940 37130 16247
rect 36793 15912 37130 15940
rect 37889 16259 38226 16286
rect 37889 15952 37918 16259
rect 38189 15952 38226 16259
rect 37889 15916 38226 15952
rect 39137 16263 39474 16286
rect 39137 15956 39169 16263
rect 39440 15956 39474 16263
rect 39137 15916 39474 15956
rect 40761 16255 41098 16286
rect 40761 15948 40792 16255
rect 41063 15948 41098 16255
rect 40761 15916 41098 15948
rect 41419 16247 41756 16282
rect 41419 15940 41451 16247
rect 41722 15940 41756 16247
rect 41419 15912 41756 15940
rect 42515 16259 42852 16286
rect 42515 15952 42544 16259
rect 42815 15952 42852 16259
rect 42515 15916 42852 15952
rect 43763 16263 44100 16286
rect 43763 15956 43795 16263
rect 44066 15956 44100 16263
rect 43763 15916 44100 15956
rect 45387 16255 45724 16286
rect 45387 15948 45418 16255
rect 45689 15948 45724 16255
rect 45387 15916 45724 15948
rect 46045 16247 46382 16282
rect 46045 15940 46077 16247
rect 46348 15940 46382 16247
rect 46045 15912 46382 15940
rect 47141 16259 47478 16286
rect 47141 15952 47170 16259
rect 47441 15952 47478 16259
rect 47141 15916 47478 15952
rect 48389 16263 48726 16286
rect 48389 15956 48421 16263
rect 48692 15956 48726 16263
rect 48389 15916 48726 15956
rect 50013 16255 50350 16286
rect 50013 15948 50044 16255
rect 50315 15948 50350 16255
rect 50013 15916 50350 15948
rect 50671 16247 51008 16282
rect 50671 15940 50703 16247
rect 50974 15940 51008 16247
rect 50671 15912 51008 15940
rect 51767 16259 52104 16286
rect 51767 15952 51796 16259
rect 52067 15952 52104 16259
rect 51767 15916 52104 15952
rect 53015 16263 53352 16286
rect 53015 15956 53047 16263
rect 53318 15956 53352 16263
rect 53015 15916 53352 15956
rect 54639 16255 54976 16286
rect 54639 15948 54670 16255
rect 54941 15948 54976 16255
rect 54639 15916 54976 15948
rect 55297 16247 55634 16282
rect 55297 15940 55329 16247
rect 55600 15940 55634 16247
rect 55297 15912 55634 15940
rect 56393 16259 56730 16286
rect 56393 15952 56422 16259
rect 56693 15952 56730 16259
rect 56393 15916 56730 15952
rect 57641 16263 57978 16286
rect 57641 15956 57673 16263
rect 57944 15956 57978 16263
rect 57641 15916 57978 15956
rect 59265 16255 59602 16286
rect 59265 15948 59296 16255
rect 59567 15948 59602 16255
rect 59265 15916 59602 15948
rect 59923 16247 60260 16282
rect 59923 15940 59955 16247
rect 60226 15940 60260 16247
rect 59923 15912 60260 15940
rect 61019 16259 61356 16286
rect 61019 15952 61048 16259
rect 61319 15952 61356 16259
rect 61019 15916 61356 15952
rect 61867 16263 62204 16286
rect 61867 15956 61899 16263
rect 62170 15956 62204 16263
rect 61867 15916 62204 15956
rect 64191 16255 64528 16286
rect 64191 15948 64222 16255
rect 64493 15948 64528 16255
rect 64191 15916 64528 15948
rect 64849 16247 65186 16282
rect 64849 15940 64881 16247
rect 65152 15940 65186 16247
rect 64849 15912 65186 15940
rect 65645 16259 65982 16286
rect 65645 15952 65674 16259
rect 65945 15952 65982 16259
rect 65645 15916 65982 15952
rect 67074 16263 67411 16286
rect 67074 15956 67106 16263
rect 67377 15956 67411 16263
rect 67074 15916 67411 15956
rect 68517 16255 68854 16286
rect 68517 15948 68548 16255
rect 68819 15948 68854 16255
rect 68517 15916 68854 15948
rect 69175 16247 69512 16282
rect 69175 15940 69207 16247
rect 69478 15940 69512 16247
rect 69175 15912 69512 15940
rect 70271 16259 70608 16286
rect 70271 15952 70300 16259
rect 70571 15952 70608 16259
rect 70271 15916 70608 15952
rect 71519 16263 71856 16286
rect 71519 15956 71551 16263
rect 71822 15956 71856 16263
rect 71519 15916 71856 15956
rect 73143 16255 73480 16286
rect 73143 15948 73174 16255
rect 73445 15948 73480 16255
rect 73143 15916 73480 15948
rect 73971 16247 74308 16282
rect 73971 15940 74003 16247
rect 74274 15940 74308 16247
rect 73971 15912 74308 15940
rect 74897 16259 75234 16286
rect 74897 15952 74926 16259
rect 75197 15952 75234 16259
rect 74897 15916 75234 15952
rect 76145 16263 76482 16286
rect 76145 15956 76177 16263
rect 76448 15956 76482 16263
rect 76145 15916 76482 15956
rect 77769 16255 78106 16286
rect 77769 15948 77800 16255
rect 78071 15948 78106 16255
rect 77769 15916 78106 15948
rect 78597 16247 78934 16282
rect 78597 15940 78629 16247
rect 78900 15940 78934 16247
rect 78597 15912 78934 15940
rect 79523 16259 79860 16286
rect 79523 15952 79552 16259
rect 79823 15952 79860 16259
rect 79523 15916 79860 15952
rect 80771 16263 81108 16286
rect 80771 15956 80803 16263
rect 81074 15956 81108 16263
rect 80771 15916 81108 15956
rect 82395 16255 82732 16286
rect 82395 15948 82426 16255
rect 82697 15948 82732 16255
rect 82395 15916 82732 15948
rect 83053 16247 83390 16282
rect 83053 15940 83085 16247
rect 83356 15940 83390 16247
rect 83053 15912 83390 15940
rect 84149 16259 84486 16286
rect 84149 15952 84178 16259
rect 84449 15952 84486 16259
rect 84149 15916 84486 15952
rect 85397 16263 85734 16286
rect 85397 15956 85429 16263
rect 85700 15956 85734 16263
rect 85397 15916 85734 15956
rect 86921 16255 87258 16286
rect 86921 15948 86952 16255
rect 87223 15948 87258 16255
rect 86921 15916 87258 15948
rect 87849 16247 88186 16282
rect 87849 15940 87881 16247
rect 88152 15940 88186 16247
rect 87849 15912 88186 15940
rect 88775 16259 89112 16286
rect 88775 15952 88804 16259
rect 89075 15952 89112 16259
rect 88775 15916 89112 15952
rect 90023 16263 90360 16286
rect 90023 15956 90055 16263
rect 90326 15956 90360 16263
rect 90023 15916 90360 15956
rect 91647 16255 91984 16286
rect 91647 15948 91678 16255
rect 91949 15948 91984 16255
rect 91647 15916 91984 15948
rect 92505 16247 92842 16282
rect 92505 15940 92537 16247
rect 92808 15940 92842 16247
rect 92505 15912 92842 15940
rect 93401 16259 93738 16286
rect 93401 15952 93430 16259
rect 93701 15952 93738 16259
rect 93401 15916 93738 15952
rect 94649 16263 94986 16286
rect 94649 15956 94681 16263
rect 94952 15956 94986 16263
rect 94649 15916 94986 15956
rect 96073 16255 96410 16286
rect 96073 15948 96104 16255
rect 96375 15948 96410 16255
rect 96073 15916 96410 15948
rect 97031 16247 97368 16282
rect 97031 15940 97063 16247
rect 97334 15940 97368 16247
rect 97031 15912 97368 15940
rect 98027 16259 98364 16286
rect 98027 15952 98056 16259
rect 98327 15952 98364 16259
rect 98027 15916 98364 15952
rect 98575 16263 98912 16286
rect 98575 15956 98607 16263
rect 98878 15956 98912 16263
rect 98575 15916 98912 15956
rect 100699 16255 101036 16286
rect 100699 15948 100730 16255
rect 101001 15948 101036 16255
rect 100699 15916 101036 15948
rect 101757 16247 102094 16282
rect 101757 15940 101789 16247
rect 102060 15940 102094 16247
rect 101757 15912 102094 15940
rect 102653 16259 102990 16286
rect 102653 15952 102682 16259
rect 102953 15952 102990 16259
rect 102653 15916 102990 15952
rect 103901 16263 104238 16286
rect 103901 15956 103933 16263
rect 104204 15956 104238 16263
rect 103901 15916 104238 15956
rect 105125 16255 105462 16286
rect 105125 15948 105156 16255
rect 105427 15948 105462 16255
rect 105125 15916 105462 15948
rect 106383 16247 106720 16282
rect 106383 15940 106415 16247
rect 106686 15940 106720 16247
rect 106383 15912 106720 15940
rect 107279 16259 107616 16286
rect 107279 15952 107308 16259
rect 107579 15952 107616 16259
rect 107279 15916 107616 15952
rect 108527 16263 108864 16286
rect 108527 15956 108559 16263
rect 108830 15956 108864 16263
rect 108527 15916 108864 15956
rect 110051 16255 110388 16286
rect 110051 15948 110082 16255
rect 110353 15948 110388 16255
rect 110051 15916 110388 15948
rect 111009 16247 111346 16282
rect 111009 15940 111041 16247
rect 111312 15940 111346 16247
rect 111009 15912 111346 15940
rect 111905 16259 112242 16286
rect 111905 15952 111934 16259
rect 112205 15952 112242 16259
rect 111905 15916 112242 15952
rect 113153 16263 113490 16286
rect 113153 15956 113185 16263
rect 113456 15956 113490 16263
rect 113153 15916 113490 15956
rect 114777 16255 115114 16286
rect 114777 15948 114808 16255
rect 115079 15948 115114 16255
rect 114777 15916 115114 15948
rect 115635 16247 115972 16282
rect 115635 15940 115667 16247
rect 115938 15940 115972 16247
rect 115635 15912 115972 15940
rect 116531 16259 116868 16286
rect 116531 15952 116560 16259
rect 116831 15952 116868 16259
rect 116531 15916 116868 15952
rect 117779 16263 118116 16286
rect 117779 15956 117811 16263
rect 118082 15956 118116 16263
rect 117779 15916 118116 15956
rect 119303 16255 119640 16286
rect 119303 15948 119334 16255
rect 119605 15948 119640 16255
rect 119303 15916 119640 15948
rect 120261 16247 120598 16282
rect 120261 15940 120293 16247
rect 120564 15940 120598 16247
rect 120261 15912 120598 15940
rect 121157 16259 121494 16286
rect 121157 15952 121186 16259
rect 121457 15952 121494 16259
rect 121157 15916 121494 15952
rect 122405 16263 122742 16286
rect 122405 15956 122437 16263
rect 122708 15956 122742 16263
rect 122405 15916 122742 15956
rect 124029 16255 124366 16286
rect 124029 15948 124060 16255
rect 124331 15948 124366 16255
rect 124029 15916 124366 15948
rect 124887 16247 125224 16282
rect 124887 15940 124919 16247
rect 125190 15940 125224 16247
rect 124887 15912 125224 15940
rect 125783 16259 126120 16286
rect 125783 15952 125812 16259
rect 126083 15952 126120 16259
rect 125783 15916 126120 15952
rect 127031 16263 127368 16286
rect 127031 15956 127063 16263
rect 127334 15956 127368 16263
rect 127031 15916 127368 15956
rect 128455 16255 128792 16286
rect 128455 15948 128486 16255
rect 128757 15948 128792 16255
rect 128455 15916 128792 15948
rect 129513 16247 129850 16282
rect 129513 15940 129545 16247
rect 129816 15940 129850 16247
rect 129513 15912 129850 15940
rect 130409 16259 130746 16286
rect 130409 15952 130438 16259
rect 130709 15952 130746 16259
rect 130409 15916 130746 15952
rect 131657 16263 131994 16286
rect 131657 15956 131689 16263
rect 131960 15956 131994 16263
rect 131657 15916 131994 15956
rect 133281 16255 133618 16286
rect 133281 15948 133312 16255
rect 133583 15948 133618 16255
rect 133281 15916 133618 15948
rect 133839 16247 134176 16282
rect 133839 15940 133871 16247
rect 134142 15940 134176 16247
rect 133839 15912 134176 15940
rect 135035 16259 135372 16286
rect 135035 15952 135064 16259
rect 135335 15952 135372 16259
rect 135035 15916 135372 15952
rect 136283 16263 136620 16286
rect 136283 15956 136315 16263
rect 136586 15956 136620 16263
rect 136283 15916 136620 15956
rect 137907 16255 138244 16286
rect 137907 15948 137938 16255
rect 138209 15948 138244 16255
rect 137907 15916 138244 15948
use cv3_via2_6cut  cv3_via2_6cut_0
timestamp 1719259570
transform 1 0 9344 0 1 2
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_1
timestamp 1719259570
transform 1 0 37100 0 1 514
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_2
timestamp 1719259570
transform 1 0 92 0 1 2
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_3
timestamp 1719259570
transform 1 0 4718 0 1 2
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_4
timestamp 1719259570
transform 1 0 13970 0 1 2
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_5
timestamp 1719259570
transform 1 0 36539 0 1 7684
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_6
timestamp 1719259570
transform 1 0 50978 0 1 1026
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_7
timestamp 1719259570
transform 1 0 129621 0 1 7170
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_8
timestamp 1719259570
transform 1 0 23208 0 1 515
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_9
timestamp 1719259570
transform 1 0 69482 0 1 1538
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_10
timestamp 1719259570
transform 1 0 41726 0 1 514
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_11
timestamp 1719259570
transform 1 0 46352 0 1 1026
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_12
timestamp 1719259570
transform 1 0 50397 0 1 5114
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_13
timestamp 1719259570
transform 1 0 74108 0 1 1538
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_14
timestamp 1719259570
transform 1 0 78734 0 1 1538
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_15
timestamp 1719259570
transform 1 0 64856 0 1 1026
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_16
timestamp 1719259570
transform 1 0 22654 0 1 3579
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_17
timestamp 1719259570
transform 1 0 83360 0 1 1538
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_18
timestamp 1719259570
transform 1 0 22684 0 1 12804
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_19
timestamp 1719259570
transform 1 0 96669 0 1 10237
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_20
timestamp 1719259570
transform 1 0 13405 0 1 8190
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_21
timestamp 1719259570
transform 1 0 18596 0 1 2
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_22
timestamp 1719259570
transform 1 0 32474 0 1 514
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_23
timestamp 1719259570
transform 1 0 27849 0 1 509
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_24
timestamp 1719259570
transform 1 0 101295 0 1 6149
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_25
timestamp 1719259570
transform 1 0 97238 0 1 2050
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_26
timestamp 1719259570
transform 1 0 101864 0 1 2050
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_27
timestamp 1719259570
transform 1 0 111122 0 1 6667
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_28
timestamp 1719259570
transform 1 0 27277 0 1 10751
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_29
timestamp 1719259570
transform 1 0 31899 0 1 11796
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_30
timestamp 1719259570
transform 1 0 87986 0 1 1538
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_31
timestamp 1719259570
transform 1 0 -484 0 1 4090
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_32
timestamp 1719259570
transform 1 0 -477 0 1 13309
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_33
timestamp 1719259570
transform 1 0 50397 0 1 11264
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_34
timestamp 1719259570
transform 1 0 8817 0 1 12301
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_35
timestamp 1719259570
transform 1 0 45788 0 1 4102
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_36
timestamp 1719259570
transform 1 0 8778 0 1 6138
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_37
timestamp 1719259570
transform 1 0 13386 0 1 9216
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_38
timestamp 1719259570
transform 1 0 60230 0 1 1026
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_39
timestamp 1719259570
transform 1 0 55604 0 1 1026
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_40
timestamp 1719259570
transform 1 0 45803 0 1 13296
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_41
timestamp 1719259570
transform 1 0 41151 0 1 9720
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_42
timestamp 1719259570
transform 1 0 4137 0 1 5114
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_43
timestamp 1719259570
transform 1 0 55038 0 1 6138
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_44
timestamp 1719259570
transform 1 0 59665 0 1 8190
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_45
timestamp 1719259570
transform 1 0 59646 0 1 9216
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_46
timestamp 1719259570
transform 1 0 4137 0 1 11264
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_47
timestamp 1719259570
transform 1 0 64287 0 1 10251
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_48
timestamp 1719259570
transform 1 0 55077 0 1 12301
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_49
timestamp 1719259570
transform 1 0 82800 0 1 8710
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_50
timestamp 1719259570
transform 1 0 92049 0 1 8198
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_51
timestamp 1719259570
transform 1 0 78159 0 1 11796
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_52
timestamp 1719259570
transform 1 0 73537 0 1 10751
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_53
timestamp 1719259570
transform 1 0 68944 0 1 12804
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_54
timestamp 1719259570
transform 1 0 18027 0 1 10251
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_55
timestamp 1719259570
transform 1 0 27271 0 1 4602
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_56
timestamp 1719259570
transform 1 0 31912 0 1 5625
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_57
timestamp 1719259570
transform 1 0 68914 0 1 3579
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_58
timestamp 1719259570
transform 1 0 73531 0 1 4602
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_59
timestamp 1719259570
transform 1 0 78172 0 1 5625
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_60
timestamp 1719259570
transform 1 0 36540 0 1 8710
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_61
timestamp 1719259570
transform 1 0 82799 0 1 7684
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_62
timestamp 1719259570
transform 1 0 87411 0 1 9720
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_63
timestamp 1719259570
transform 1 0 101292 0 1 12305
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_64
timestamp 1719259570
transform 1 0 110560 0 1 8709
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_65
timestamp 1719259570
transform 1 0 92612 0 1 2050
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_66
timestamp 1719259570
transform 1 0 92045 0 1 4108
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_67
timestamp 1719259570
transform 1 0 96675 0 1 5114
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_68
timestamp 1719259570
transform 1 0 106490 0 1 2050
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_69
timestamp 1719259570
transform 1 0 134247 0 1 7170
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_70
timestamp 1719259570
transform 1 0 115728 0 1 6667
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_71
timestamp 1719259570
transform 1 0 120375 0 1 6667
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_72
timestamp 1719259570
transform 1 0 124984 0 1 7170
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_73
timestamp 1719259570
transform 1 0 105921 0 1 13310
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_74
timestamp 1719259570
transform 1 0 110556 0 1 3588
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_75
timestamp 1719259570
transform 1 0 115168 0 1 10758
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_76
timestamp 1719259570
transform 1 0 124434 0 1 4087
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_77
timestamp 1719259570
transform 1 0 119794 0 1 5621
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_78
timestamp 1719259570
transform 1 0 133684 0 1 6150
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_79
timestamp 1719259570
transform 1 0 129050 0 1 5126
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_80
timestamp 1719259570
transform 1 0 129054 0 1 11776
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_81
timestamp 1719259570
transform 1 0 124428 0 1 9726
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_82
timestamp 1719259570
transform 1 0 115156 0 1 4618
box 3030 432 3561 574
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_0 ../dependencies/sky130_ef_ip__analog_switches/mag
array 0 0 -3542 0 29 -4626
timestamp 1724439637
transform 0 -1 3580 -1 0 7619
box -4 -600 3538 3648
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_1
array 0 0 -3542 0 3 -4626
timestamp 1724439637
transform 0 -1 49843 -1 0 13272
box -4 -600 3538 3648
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_2
array 0 0 -3542 0 3 -4626
timestamp 1724439637
transform 0 -1 3583 -1 0 13272
box -4 -600 3538 3648
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_3
array 0 0 -3542 0 3 -4626
timestamp 1724439637
transform 0 -1 26713 -1 0 13272
box -4 -600 3538 3648
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_4
array 0 0 -3542 0 1 -4626
timestamp 1724439637
transform 0 -1 128485 -1 0 13272
box -4 -600 3538 3648
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_5
array 0 0 -3542 0 3 -4626
timestamp 1724439637
transform 0 -1 72973 -1 0 13272
box -4 -600 3538 3648
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_6
array 0 0 -3542 0 2 -4626
timestamp 1724439637
transform 0 -1 96103 -1 0 13272
box -4 -600 3538 3648
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_7
array 0 0 -3542 0 1 -4626
timestamp 1724439637
transform 0 -1 114607 -1 0 13272
box -4 -600 3538 3648
<< labels >>
flabel comment s -843 13866 -843 13866 0 FreeSans 960 0 0 0 right_instramp_p
flabel comment s -425 13354 -425 13354 0 FreeSans 960 0 0 0 right_instramp_n
flabel comment s -449 12838 -449 12838 0 FreeSans 960 0 0 0 right_lp_opamp_p
flabel comment s -517 12324 -517 12324 0 FreeSans 960 0 0 0 right_lp_opamp_n
flabel comment s -527 11820 -527 11820 0 FreeSans 960 0 0 0 right_hgbw_opamp_p
flabel comment s -449 11302 -449 11302 0 FreeSans 960 0 0 0 right_hgbw_opamp_n
flabel comment s -455 10794 -455 10794 0 FreeSans 960 0 0 0 left_hgbw_opamp_p
flabel comment s -471 10288 -471 10288 0 FreeSans 960 0 0 0 left_hgbw_opamp_n
flabel comment s -479 9768 -479 9768 0 FreeSans 960 0 0 0 left_lp_opamp_p
flabel comment s -519 9266 -519 9266 0 FreeSans 960 0 0 0 left_lp_opamp_n
flabel comment s -477 8748 -477 8748 0 FreeSans 960 0 0 0 left_instramp_p
flabel comment s -493 8232 -493 8232 0 FreeSans 960 0 0 0 left_instramp_n
flabel comment s -553 7722 -553 7722 0 FreeSans 960 0 0 0 vbgtc
flabel comment s -567 7204 -567 7204 0 FreeSans 960 0 0 0 vbgsc
flabel comment s -579 6702 -579 6702 0 FreeSans 960 0 0 0 ulp_comp_p
flabel comment s -607 6184 -607 6184 0 FreeSans 960 0 0 0 ulp_comp_n
flabel comment s -643 5672 -643 5672 0 FreeSans 960 0 0 0 comp_p
flabel comment s -681 5160 -681 5160 0 FreeSans 960 0 0 0 comp_n
flabel comment s -689 4648 -689 4648 0 FreeSans 960 0 0 0 adc0_in
flabel comment s -679 4136 -679 4136 0 FreeSans 960 0 0 0 adc1_in
flabel comment s -675 2600 -675 2600 0 FreeSans 960 0 0 0 tempsense_out
flabel comment s -659 2086 -659 2086 0 FreeSans 960 0 0 0 right_vref
flabel comment s -667 1578 -667 1578 0 FreeSans 960 0 0 0 left_vref
flabel comment s -663 1074 -663 1074 0 FreeSans 960 0 0 0 vinref
flabel comment s -689 554 -689 554 0 FreeSans 960 0 0 0 voutref
flabel comment s 139384 525 139384 525 0 FreeSans 960 0 0 0 voutref
flabel comment s 139410 1045 139410 1045 0 FreeSans 960 0 0 0 vinref
flabel comment s 139406 1549 139406 1549 0 FreeSans 960 0 0 0 left_vref
flabel comment s 139414 2057 139414 2057 0 FreeSans 960 0 0 0 right_vref
flabel comment s 139398 2571 139398 2571 0 FreeSans 960 0 0 0 tempsense_out
flabel comment s 139394 4107 139394 4107 0 FreeSans 960 0 0 0 adc1_in
flabel comment s 139384 4619 139384 4619 0 FreeSans 960 0 0 0 adc0_in
flabel comment s 139392 5131 139392 5131 0 FreeSans 960 0 0 0 comp_n
flabel comment s 139430 5643 139430 5643 0 FreeSans 960 0 0 0 comp_p
flabel comment s 139466 6155 139466 6155 0 FreeSans 960 0 0 0 ulp_comp_n
flabel comment s 139494 6673 139494 6673 0 FreeSans 960 0 0 0 ulp_comp_p
flabel comment s 139506 7175 139506 7175 0 FreeSans 960 0 0 0 vbgsc
flabel comment s 139520 7693 139520 7693 0 FreeSans 960 0 0 0 vbgtc
flabel comment s 139580 8203 139580 8203 0 FreeSans 960 0 0 0 left_instramp_n
flabel comment s 139596 8719 139596 8719 0 FreeSans 960 0 0 0 left_instramp_p
flabel comment s 139554 9237 139554 9237 0 FreeSans 960 0 0 0 left_lp_opamp_n
flabel comment s 139594 9739 139594 9739 0 FreeSans 960 0 0 0 left_lp_opamp_p
flabel comment s 139602 10259 139602 10259 0 FreeSans 960 0 0 0 left_hgbw_opamp_n
flabel comment s 139618 10765 139618 10765 0 FreeSans 960 0 0 0 left_hgbw_opamp_p
flabel comment s 139624 11273 139624 11273 0 FreeSans 960 0 0 0 right_hgbw_opamp_n
flabel comment s 139546 11791 139546 11791 0 FreeSans 960 0 0 0 right_hgbw_opamp_p
flabel comment s 139556 12295 139556 12295 0 FreeSans 960 0 0 0 right_lp_opamp_n
flabel comment s 139624 12809 139624 12809 0 FreeSans 960 0 0 0 right_lp_opamp_p
flabel comment s 139648 13325 139648 13325 0 FreeSans 960 0 0 0 right_instramp_n
flabel comment s 139230 13837 139230 13837 0 FreeSans 960 0 0 0 right_instramp_p
<< end >>
