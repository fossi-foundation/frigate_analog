magic
tech sky130A
magscale 1 2
timestamp 1716557812
<< checkpaint >>
rect 166206 106631 185634 107641
rect 166108 106325 189814 106631
rect 166108 106249 190120 106325
rect 194862 106249 214290 107641
rect 103854 103703 165438 104107
rect 166108 103703 214290 106249
rect 279926 104107 301766 116578
rect 345662 114349 504708 127977
rect 223782 103703 301766 104107
rect 103854 78452 301766 103703
rect 330502 105303 504708 114349
rect 330502 85614 512236 105303
rect 108134 78048 268938 78452
rect 108134 77972 207688 78048
rect 170692 77666 207688 77972
rect 188260 77590 207688 77666
rect 279926 63958 301766 78452
rect 330656 79648 512236 85614
rect 330656 77346 489854 79648
rect 330656 77040 489702 77346
rect 20584 55468 30298 57444
rect 20584 51334 38930 55468
rect 14398 50764 38930 51334
rect 279926 52450 349822 63958
rect 12118 8814 39174 50764
rect 262580 48770 275674 50480
rect 12118 8244 25212 8814
rect 26080 8244 39174 8814
rect 260586 7960 275674 48770
rect 279926 8330 351296 52450
rect 471410 34760 516553 58771
rect 564880 56488 618644 64026
rect 528546 26232 556148 50338
rect 260586 6250 273680 7960
rect 10622 -5218 13376 516
rect 279926 -1260 301766 8330
rect 412740 -54726 425834 -12206
<< comment >>
rect 58 109226 627978 115318
rect 0 105318 627978 109226
rect 0 78620 10124 105318
rect 20160 80752 96352 100466
rect 281186 78620 294506 105318
rect 515230 82052 591422 101766
rect 618596 78620 627978 105318
rect 0 58620 627978 78620
rect 0 4758 10124 58620
rect 46166 7586 83464 54474
rect 93052 7052 130350 53940
rect 136210 7586 173508 54474
rect 178302 8118 215600 55006
rect 219330 7052 256628 53940
rect 281186 4758 294506 58620
rect 347386 4758 362304 58620
rect 371104 22910 418790 55944
rect 529806 27492 554888 49078
rect 566912 24508 614866 57008
rect 618596 4758 627978 58620
rect 0 0 627978 4758
use bias_generator  bias_generator_0 ../ip/sky130_ef_ip__biasgen/mag
timestamp 1715390562
transform 1 0 367174 0 1 15943
box -1132 -6353 249191 3114
use sky130_ak_ip__comparator  sky130_ak_ip__comparator_0 ../ip/sky130_ak_ip__comparator/mag
timestamp 1715629873
transform 0 1 331006 -1 0 55784
box -1900 -33700 39700 13700
use sky130_cw_ip__bandgap  sky130_cw_ip__bandgap_0 ../ip/sky130_cw_ip/mag
timestamp 1715625863
transform 1 0 427432 0 1 43290
box -5734 12 42048 14837
use sky130_ef_ip__rheostat_8bit  sky130_ef_ip__rheostat_8bit_0 ../ip/sky130_ef_ip__rheostat_8bit/mag
timestamp 1716082924
transform 0 1 189524 1 0 79050
box -200 -4 25939 16904
use sky130_ef_ip__rheostat_8bit  sky130_ef_ip__rheostat_8bit_1
timestamp 1716082924
transform 0 -1 188856 1 0 79126
box -200 -4 25939 16904
use sky130_ef_ip__rheostat_8bit  sky130_ef_ip__rheostat_8bit_2
timestamp 1716082924
transform 0 1 410440 1 0 79112
box -200 -4 25939 16904
use sky130_ef_ip__rheostat_8bit  sky130_ef_ip__rheostat_8bit_3
timestamp 1716082924
transform 0 -1 409772 1 0 79188
box -200 -4 25939 16904
use sky130_fd_io__top_pwrdetv2  sky130_fd_io__top_pwrdetv2_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1715205430
transform 1 0 27058 0 1 9504
box 282 0 10856 40000
use sky130_fd_io__top_pwrdetv2  sky130_fd_io__top_pwrdetv2_1
timestamp 1715205430
transform 1 0 13096 0 1 9504
box 282 0 10856 40000
use sky130_od_ip__tempsensor_ext_vp  sky130_od_ip__tempsensor_ext_vp_0 ../ip/sky130_od_ip__tempsensor/mag
timestamp 1715712088
transform 1 0 264424 0 1 13680
box -584 -5030 6610 3202
use sky130_td_ip__opamp_hp  sky130_td_ip__opamp_hp_0 ../ip/sky130_td_ip__opamp_hp/mag
timestamp 1714591961
transform 1 0 437254 0 1 86299
box -7724 -6929 51340 16206
use sky130_td_ip__opamp_hp  sky130_td_ip__opamp_hp_1
timestamp 1714591961
transform -1 0 383408 0 1 86299
box -7724 -6929 51340 16206
use sky130_td_ip__opamp_hp  sky130_td_ip__opamp_hp_2
timestamp 1714591961
transform 1 0 216338 0 1 86237
box -7724 -6929 51340 16206
use sky130_td_ip__opamp_hp  sky130_td_ip__opamp_hp_3
timestamp 1714591961
transform -1 0 162492 0 1 86237
box -7724 -6929 51340 16206
use sky130_vbl_ip__overvoltage  sky130_vbl_ip__overvoltage_0 ../ip/sky130_vbl_ip__overvoltage/mag
timestamp 1714660490
transform 1 0 490888 0 1 40022
box -18218 -4002 24405 17489
<< labels >>
flabel comment 553592 90844 553592 90844 0 FreeSans 80000 0 0 0 inst_amp
flabel comment 371104 22910 399608 55944 0 FreeSans 80000 0 0 0 ULP_comp
flabel comment 591422 39162 591422 39162 0 FreeSans 80000 0 0 0 iDAC
flabel comment 111168 29698 111168 29698 0 FreeSans 80000 0 0 0 RDAC
flabel comment 155126 30762 155126 30762 0 FreeSans 80000 0 0 0 RDAC
flabel comment 197218 29698 197218 29698 0 FreeSans 80000 0 0 0 ADC
flabel comment 237446 28898 237446 28898 0 FreeSans 80000 0 0 0 ADC
flabel comment 64280 31030 64280 31030 0 FreeSans 80000 0 0 0 SD_DAC
flabel comment 55592 89544 55592 89544 0 FreeSans 80000 0 0 0 inst_amp
flabel comment 542750 39628 542750 39628 0 FreeSans 80000 0 0 0 POR
<< properties >>
string FIXED_BBOX 0 0 627978 115318
<< end >>
