magic
tech sky130A
magscale 1 2
timestamp 1563083296
<< checkpaint >>
rect -1260 -1260 45420 801494
<< metal2 >>
rect 19639 889 19907 941
rect 19639 433 19665 889
rect 19881 433 19907 889
rect 19639 386 19907 433
<< via2 >>
rect 19665 433 19881 889
<< metal3 >>
rect 43152 772543 43918 772575
rect 43152 772479 43185 772543
rect 43249 772479 43265 772543
rect 43329 772479 43345 772543
rect 43409 772479 43425 772543
rect 43489 772479 43505 772543
rect 43569 772479 43585 772543
rect 43649 772479 43665 772543
rect 43729 772479 43745 772543
rect 43809 772479 43825 772543
rect 43889 772479 43918 772543
rect 43152 772446 43918 772479
rect 43152 751543 43918 751575
rect 43152 751479 43185 751543
rect 43249 751479 43265 751543
rect 43329 751479 43345 751543
rect 43409 751479 43425 751543
rect 43489 751479 43505 751543
rect 43569 751479 43585 751543
rect 43649 751479 43665 751543
rect 43729 751479 43745 751543
rect 43809 751479 43825 751543
rect 43889 751479 43918 751543
rect 43152 751446 43918 751479
rect 43152 730543 43918 730575
rect 43152 730479 43185 730543
rect 43249 730479 43265 730543
rect 43329 730479 43345 730543
rect 43409 730479 43425 730543
rect 43489 730479 43505 730543
rect 43569 730479 43585 730543
rect 43649 730479 43665 730543
rect 43729 730479 43745 730543
rect 43809 730479 43825 730543
rect 43889 730479 43918 730543
rect 43152 730446 43918 730479
rect 43152 709543 43918 709575
rect 43152 709479 43185 709543
rect 43249 709479 43265 709543
rect 43329 709479 43345 709543
rect 43409 709479 43425 709543
rect 43489 709479 43505 709543
rect 43569 709479 43585 709543
rect 43649 709479 43665 709543
rect 43729 709479 43745 709543
rect 43809 709479 43825 709543
rect 43889 709479 43918 709543
rect 43152 709446 43918 709479
rect 43152 619344 43918 619353
rect 43152 619321 44160 619344
rect 43152 619257 43185 619321
rect 43249 619257 43265 619321
rect 43329 619257 43345 619321
rect 43409 619257 43425 619321
rect 43489 619257 43505 619321
rect 43569 619257 43585 619321
rect 43649 619257 43665 619321
rect 43729 619257 43745 619321
rect 43809 619257 43825 619321
rect 43889 619257 44160 619321
rect 43152 619224 44160 619257
rect 43152 586344 43918 586353
rect 43152 586321 44160 586344
rect 43152 586257 43185 586321
rect 43249 586257 43265 586321
rect 43329 586257 43345 586321
rect 43409 586257 43425 586321
rect 43489 586257 43505 586321
rect 43569 586257 43585 586321
rect 43649 586257 43665 586321
rect 43729 586257 43745 586321
rect 43809 586257 43825 586321
rect 43889 586257 44160 586321
rect 43152 586224 44160 586257
rect 43152 553344 43918 553353
rect 43152 553321 44160 553344
rect 43152 553257 43185 553321
rect 43249 553257 43265 553321
rect 43329 553257 43345 553321
rect 43409 553257 43425 553321
rect 43489 553257 43505 553321
rect 43569 553257 43585 553321
rect 43649 553257 43665 553321
rect 43729 553257 43745 553321
rect 43809 553257 43825 553321
rect 43889 553257 44160 553321
rect 43152 553224 44160 553257
rect 43152 520344 43918 520353
rect 43152 520321 44160 520344
rect 43152 520257 43185 520321
rect 43249 520257 43265 520321
rect 43329 520257 43345 520321
rect 43409 520257 43425 520321
rect 43489 520257 43505 520321
rect 43569 520257 43585 520321
rect 43649 520257 43665 520321
rect 43729 520257 43745 520321
rect 43809 520257 43825 520321
rect 43889 520257 44160 520321
rect 43152 520224 44160 520257
rect 43101 465624 43895 466024
rect 43152 456559 43918 456568
rect 43152 456536 44160 456559
rect 43152 456472 43185 456536
rect 43249 456472 43265 456536
rect 43329 456472 43345 456536
rect 43409 456472 43425 456536
rect 43489 456472 43505 456536
rect 43569 456472 43585 456536
rect 43649 456472 43665 456536
rect 43729 456472 43745 456536
rect 43809 456472 43825 456536
rect 43889 456472 44160 456536
rect 43152 456439 44160 456472
rect 43152 422744 43918 422753
rect 43152 422721 44160 422744
rect 43152 422657 43185 422721
rect 43249 422657 43265 422721
rect 43329 422657 43345 422721
rect 43409 422657 43425 422721
rect 43489 422657 43505 422721
rect 43569 422657 43585 422721
rect 43649 422657 43665 422721
rect 43729 422657 43745 422721
rect 43809 422657 43825 422721
rect 43889 422657 44160 422721
rect 43152 422624 44160 422657
rect 43152 389744 43918 389753
rect 43152 389721 44160 389744
rect 43152 389657 43185 389721
rect 43249 389657 43265 389721
rect 43329 389657 43345 389721
rect 43409 389657 43425 389721
rect 43489 389657 43505 389721
rect 43569 389657 43585 389721
rect 43649 389657 43665 389721
rect 43729 389657 43745 389721
rect 43809 389657 43825 389721
rect 43889 389657 44160 389721
rect 43152 389624 44160 389657
rect 43152 356487 43918 356496
rect 43152 356464 44160 356487
rect 43152 356400 43185 356464
rect 43249 356400 43265 356464
rect 43329 356400 43345 356464
rect 43409 356400 43425 356464
rect 43489 356400 43505 356464
rect 43569 356400 43585 356464
rect 43649 356400 43665 356464
rect 43729 356400 43745 356464
rect 43809 356400 43825 356464
rect 43889 356400 44160 356464
rect 43152 356367 44160 356400
rect 43152 323487 43918 323496
rect 43152 323464 44160 323487
rect 43152 323400 43185 323464
rect 43249 323400 43265 323464
rect 43329 323400 43345 323464
rect 43409 323400 43425 323464
rect 43489 323400 43505 323464
rect 43569 323400 43585 323464
rect 43649 323400 43665 323464
rect 43729 323400 43745 323464
rect 43809 323400 43825 323464
rect 43889 323400 44160 323464
rect 43152 323367 44160 323400
rect 19531 962 19906 1000
rect 19531 418 19564 962
rect 19868 889 19906 962
rect 19881 433 19906 889
rect 19868 418 19906 433
rect 19531 386 19906 418
<< via3 >>
rect 43185 772479 43249 772543
rect 43265 772479 43329 772543
rect 43345 772479 43409 772543
rect 43425 772479 43489 772543
rect 43505 772479 43569 772543
rect 43585 772479 43649 772543
rect 43665 772479 43729 772543
rect 43745 772479 43809 772543
rect 43825 772479 43889 772543
rect 43185 751479 43249 751543
rect 43265 751479 43329 751543
rect 43345 751479 43409 751543
rect 43425 751479 43489 751543
rect 43505 751479 43569 751543
rect 43585 751479 43649 751543
rect 43665 751479 43729 751543
rect 43745 751479 43809 751543
rect 43825 751479 43889 751543
rect 43185 730479 43249 730543
rect 43265 730479 43329 730543
rect 43345 730479 43409 730543
rect 43425 730479 43489 730543
rect 43505 730479 43569 730543
rect 43585 730479 43649 730543
rect 43665 730479 43729 730543
rect 43745 730479 43809 730543
rect 43825 730479 43889 730543
rect 43185 709479 43249 709543
rect 43265 709479 43329 709543
rect 43345 709479 43409 709543
rect 43425 709479 43489 709543
rect 43505 709479 43569 709543
rect 43585 709479 43649 709543
rect 43665 709479 43729 709543
rect 43745 709479 43809 709543
rect 43825 709479 43889 709543
rect 43185 619257 43249 619321
rect 43265 619257 43329 619321
rect 43345 619257 43409 619321
rect 43425 619257 43489 619321
rect 43505 619257 43569 619321
rect 43585 619257 43649 619321
rect 43665 619257 43729 619321
rect 43745 619257 43809 619321
rect 43825 619257 43889 619321
rect 43185 586257 43249 586321
rect 43265 586257 43329 586321
rect 43345 586257 43409 586321
rect 43425 586257 43489 586321
rect 43505 586257 43569 586321
rect 43585 586257 43649 586321
rect 43665 586257 43729 586321
rect 43745 586257 43809 586321
rect 43825 586257 43889 586321
rect 43185 553257 43249 553321
rect 43265 553257 43329 553321
rect 43345 553257 43409 553321
rect 43425 553257 43489 553321
rect 43505 553257 43569 553321
rect 43585 553257 43649 553321
rect 43665 553257 43729 553321
rect 43745 553257 43809 553321
rect 43825 553257 43889 553321
rect 43185 520257 43249 520321
rect 43265 520257 43329 520321
rect 43345 520257 43409 520321
rect 43425 520257 43489 520321
rect 43505 520257 43569 520321
rect 43585 520257 43649 520321
rect 43665 520257 43729 520321
rect 43745 520257 43809 520321
rect 43825 520257 43889 520321
rect 43185 456472 43249 456536
rect 43265 456472 43329 456536
rect 43345 456472 43409 456536
rect 43425 456472 43489 456536
rect 43505 456472 43569 456536
rect 43585 456472 43649 456536
rect 43665 456472 43729 456536
rect 43745 456472 43809 456536
rect 43825 456472 43889 456536
rect 43185 422657 43249 422721
rect 43265 422657 43329 422721
rect 43345 422657 43409 422721
rect 43425 422657 43489 422721
rect 43505 422657 43569 422721
rect 43585 422657 43649 422721
rect 43665 422657 43729 422721
rect 43745 422657 43809 422721
rect 43825 422657 43889 422721
rect 43185 389657 43249 389721
rect 43265 389657 43329 389721
rect 43345 389657 43409 389721
rect 43425 389657 43489 389721
rect 43505 389657 43569 389721
rect 43585 389657 43649 389721
rect 43665 389657 43729 389721
rect 43745 389657 43809 389721
rect 43825 389657 43889 389721
rect 43185 356400 43249 356464
rect 43265 356400 43329 356464
rect 43345 356400 43409 356464
rect 43425 356400 43489 356464
rect 43505 356400 43569 356464
rect 43585 356400 43649 356464
rect 43665 356400 43729 356464
rect 43745 356400 43809 356464
rect 43825 356400 43889 356464
rect 43185 323400 43249 323464
rect 43265 323400 43329 323464
rect 43345 323400 43409 323464
rect 43425 323400 43489 323464
rect 43505 323400 43569 323464
rect 43585 323400 43649 323464
rect 43665 323400 43729 323464
rect 43745 323400 43809 323464
rect 43825 323400 43889 323464
rect 19564 889 19868 962
rect 19564 433 19665 889
rect 19665 433 19868 889
rect 19564 418 19868 433
<< metal4 >>
rect 535 317481 663 800234
rect 795 317741 923 800234
rect 1047 317993 1175 800234
rect 1307 318253 1435 800234
rect 1559 318505 1687 800234
rect 1819 318765 1947 800234
rect 2071 319017 2199 800234
rect 2331 319277 2459 800234
rect 2583 319529 2711 800234
rect 2843 319789 2971 800234
rect 3095 320041 3223 800234
rect 3355 320301 3483 800234
rect 3607 320553 3735 800234
rect 3867 320813 3995 800234
rect 4119 321065 4247 800234
rect 4379 323597 4507 800234
rect 4639 324284 4767 800234
rect 4891 356568 5019 800234
rect 5151 357268 5279 800234
rect 5403 389853 5531 800234
rect 5663 390487 5791 800234
rect 5915 422854 6043 800234
rect 6175 423449 6303 800234
rect 6427 456669 6555 800234
rect 6687 457224 6815 800234
rect 6939 520454 7067 800234
rect 7199 521024 7327 800234
rect 7451 553454 7579 800234
rect 7711 554144 7839 800234
rect 7963 586454 8091 800234
rect 8223 587083 8351 800234
rect 8475 619435 8603 800234
rect 8735 620146 8863 800234
rect 8987 709676 9115 800234
rect 9247 710319 9375 800234
rect 9499 730682 9627 800234
rect 9759 731297 9887 800234
rect 10011 751692 10139 800234
rect 10271 752366 10399 800234
rect 10523 772676 10651 800234
rect 10783 773425 10911 800234
rect 42892 772635 43581 772676
rect 42892 772399 42960 772635
rect 43196 772543 43280 772635
rect 43516 772575 43581 772635
rect 43516 772543 43918 772575
rect 43249 772479 43265 772543
rect 43569 772479 43585 772543
rect 43649 772479 43665 772543
rect 43729 772479 43745 772543
rect 43809 772479 43825 772543
rect 43889 772479 43918 772543
rect 43196 772399 43280 772479
rect 43516 772446 43918 772479
rect 43516 772399 43581 772446
rect 42892 772356 43581 772399
rect 42892 751635 43581 751676
rect 42892 751399 42960 751635
rect 43196 751543 43280 751635
rect 43516 751575 43581 751635
rect 43516 751543 43918 751575
rect 43249 751479 43265 751543
rect 43569 751479 43585 751543
rect 43649 751479 43665 751543
rect 43729 751479 43745 751543
rect 43809 751479 43825 751543
rect 43889 751479 43918 751543
rect 43196 751399 43280 751479
rect 43516 751446 43918 751479
rect 43516 751399 43581 751446
rect 42892 751356 43581 751399
rect 42892 730635 43581 730676
rect 42892 730399 42960 730635
rect 43196 730543 43280 730635
rect 43516 730575 43581 730635
rect 43516 730543 43918 730575
rect 43249 730479 43265 730543
rect 43569 730479 43585 730543
rect 43649 730479 43665 730543
rect 43729 730479 43745 730543
rect 43809 730479 43825 730543
rect 43889 730479 43918 730543
rect 43196 730399 43280 730479
rect 43516 730446 43918 730479
rect 43516 730399 43581 730446
rect 42892 730356 43581 730399
rect 42892 709635 43581 709676
rect 42892 709399 42960 709635
rect 43196 709543 43280 709635
rect 43516 709575 43581 709635
rect 43516 709543 43918 709575
rect 43249 709479 43265 709543
rect 43569 709479 43585 709543
rect 43649 709479 43665 709543
rect 43729 709479 43745 709543
rect 43809 709479 43825 709543
rect 43889 709479 43918 709543
rect 43196 709399 43280 709479
rect 43516 709446 43918 709479
rect 43516 709399 43581 709446
rect 42892 709356 43581 709399
rect 42892 619413 43581 619454
rect 42892 619177 42960 619413
rect 43196 619321 43280 619413
rect 43516 619353 43581 619413
rect 43516 619321 43918 619353
rect 43249 619257 43265 619321
rect 43569 619257 43585 619321
rect 43649 619257 43665 619321
rect 43729 619257 43745 619321
rect 43809 619257 43825 619321
rect 43889 619257 43918 619321
rect 43196 619177 43280 619257
rect 43516 619224 43918 619257
rect 43516 619177 43581 619224
rect 42892 619134 43581 619177
rect 42892 586413 43581 586454
rect 42892 586177 42960 586413
rect 43196 586321 43280 586413
rect 43516 586353 43581 586413
rect 43516 586321 43918 586353
rect 43249 586257 43265 586321
rect 43569 586257 43585 586321
rect 43649 586257 43665 586321
rect 43729 586257 43745 586321
rect 43809 586257 43825 586321
rect 43889 586257 43918 586321
rect 43196 586177 43280 586257
rect 43516 586224 43918 586257
rect 43516 586177 43581 586224
rect 42892 586134 43581 586177
rect 42892 553413 43581 553454
rect 42892 553177 42960 553413
rect 43196 553321 43280 553413
rect 43516 553353 43581 553413
rect 43516 553321 43918 553353
rect 43249 553257 43265 553321
rect 43569 553257 43585 553321
rect 43649 553257 43665 553321
rect 43729 553257 43745 553321
rect 43809 553257 43825 553321
rect 43889 553257 43918 553321
rect 43196 553177 43280 553257
rect 43516 553224 43918 553257
rect 43516 553177 43581 553224
rect 42892 553134 43581 553177
rect 42892 520413 43581 520454
rect 42892 520177 42960 520413
rect 43196 520321 43280 520413
rect 43516 520353 43581 520413
rect 43516 520321 43918 520353
rect 43249 520257 43265 520321
rect 43569 520257 43585 520321
rect 43649 520257 43665 520321
rect 43729 520257 43745 520321
rect 43809 520257 43825 520321
rect 43889 520257 43918 520321
rect 43196 520177 43280 520257
rect 43516 520224 43918 520257
rect 43516 520177 43581 520224
rect 42892 520134 43581 520177
rect 43129 456669 43281 466073
rect 42892 456628 43581 456669
rect 42892 456392 42960 456628
rect 43196 456536 43280 456628
rect 43516 456568 43581 456628
rect 43516 456536 43918 456568
rect 43249 456472 43265 456536
rect 43569 456472 43585 456536
rect 43649 456472 43665 456536
rect 43729 456472 43745 456536
rect 43809 456472 43825 456536
rect 43889 456472 43918 456536
rect 43196 456392 43280 456472
rect 43516 456439 43918 456472
rect 43516 456392 43581 456439
rect 42892 456349 43581 456392
rect 42892 422813 43581 422854
rect 42892 422577 42960 422813
rect 43196 422721 43280 422813
rect 43516 422753 43581 422813
rect 43516 422721 43918 422753
rect 43249 422657 43265 422721
rect 43569 422657 43585 422721
rect 43649 422657 43665 422721
rect 43729 422657 43745 422721
rect 43809 422657 43825 422721
rect 43889 422657 43918 422721
rect 43196 422577 43280 422657
rect 43516 422624 43918 422657
rect 43516 422577 43581 422624
rect 42892 422534 43581 422577
rect 42892 389813 43581 389854
rect 42892 389577 42960 389813
rect 43196 389721 43280 389813
rect 43516 389753 43581 389813
rect 43516 389721 43918 389753
rect 43249 389657 43265 389721
rect 43569 389657 43585 389721
rect 43649 389657 43665 389721
rect 43729 389657 43745 389721
rect 43809 389657 43825 389721
rect 43889 389657 43918 389721
rect 43196 389577 43280 389657
rect 43516 389624 43918 389657
rect 43516 389577 43581 389624
rect 42892 389534 43581 389577
rect 42892 356556 43581 356597
rect 42892 356320 42960 356556
rect 43196 356464 43280 356556
rect 43516 356496 43581 356556
rect 43516 356464 43918 356496
rect 43249 356400 43265 356464
rect 43569 356400 43585 356464
rect 43649 356400 43665 356464
rect 43729 356400 43745 356464
rect 43809 356400 43825 356464
rect 43889 356400 43918 356464
rect 43196 356320 43280 356400
rect 43516 356367 43918 356400
rect 43516 356320 43581 356367
rect 42892 356277 43581 356320
rect 42892 323556 43581 323597
rect 42892 323320 42960 323556
rect 43196 323464 43280 323556
rect 43516 323496 43581 323556
rect 43516 323464 43918 323496
rect 43249 323400 43265 323464
rect 43569 323400 43585 323464
rect 43649 323400 43665 323464
rect 43729 323400 43745 323464
rect 43809 323400 43825 323464
rect 43889 323400 43918 323464
rect 43196 323320 43280 323400
rect 43516 323367 43918 323400
rect 43516 323320 43581 323367
rect 42892 323277 43581 323320
rect 4119 320937 14247 321065
rect 3867 320685 13995 320813
rect 3607 320425 13735 320553
rect 3355 320173 13483 320301
rect 3095 319913 13223 320041
rect 2843 319661 12971 319789
rect 2583 319401 12711 319529
rect 2331 319149 12459 319277
rect 2071 318889 12199 319017
rect 1819 318637 11947 318765
rect 1559 318377 11687 318505
rect 1307 318125 11435 318253
rect 1047 317865 11175 317993
rect 795 317613 10923 317741
rect 10535 317481 10663 317482
rect 535 317356 10663 317481
rect 6274 317353 10663 317356
rect 10535 12187 10663 317353
rect 10795 11180 10923 317613
rect 11047 10123 11175 317865
rect 11307 9160 11435 318125
rect 11559 8119 11687 318377
rect 11819 7285 11947 318637
rect 12071 5974 12199 318889
rect 12331 4990 12459 319149
rect 12583 4143 12711 319401
rect 12843 3304 12971 319661
rect 13095 1989 13223 319913
rect 13355 1323 13483 320173
rect 13607 0 13735 320425
rect 13867 1324 13995 320685
rect 14119 1934 14247 320937
rect 19532 962 19906 1322
rect 19532 418 19564 962
rect 19868 418 19906 962
rect 19532 387 19906 418
<< via4 >>
rect 42960 772543 43196 772635
rect 43280 772543 43516 772635
rect 42960 772479 43185 772543
rect 43185 772479 43196 772543
rect 43280 772479 43329 772543
rect 43329 772479 43345 772543
rect 43345 772479 43409 772543
rect 43409 772479 43425 772543
rect 43425 772479 43489 772543
rect 43489 772479 43505 772543
rect 43505 772479 43516 772543
rect 42960 772399 43196 772479
rect 43280 772399 43516 772479
rect 42960 751543 43196 751635
rect 43280 751543 43516 751635
rect 42960 751479 43185 751543
rect 43185 751479 43196 751543
rect 43280 751479 43329 751543
rect 43329 751479 43345 751543
rect 43345 751479 43409 751543
rect 43409 751479 43425 751543
rect 43425 751479 43489 751543
rect 43489 751479 43505 751543
rect 43505 751479 43516 751543
rect 42960 751399 43196 751479
rect 43280 751399 43516 751479
rect 42960 730543 43196 730635
rect 43280 730543 43516 730635
rect 42960 730479 43185 730543
rect 43185 730479 43196 730543
rect 43280 730479 43329 730543
rect 43329 730479 43345 730543
rect 43345 730479 43409 730543
rect 43409 730479 43425 730543
rect 43425 730479 43489 730543
rect 43489 730479 43505 730543
rect 43505 730479 43516 730543
rect 42960 730399 43196 730479
rect 43280 730399 43516 730479
rect 42960 709543 43196 709635
rect 43280 709543 43516 709635
rect 42960 709479 43185 709543
rect 43185 709479 43196 709543
rect 43280 709479 43329 709543
rect 43329 709479 43345 709543
rect 43345 709479 43409 709543
rect 43409 709479 43425 709543
rect 43425 709479 43489 709543
rect 43489 709479 43505 709543
rect 43505 709479 43516 709543
rect 42960 709399 43196 709479
rect 43280 709399 43516 709479
rect 42960 619321 43196 619413
rect 43280 619321 43516 619413
rect 42960 619257 43185 619321
rect 43185 619257 43196 619321
rect 43280 619257 43329 619321
rect 43329 619257 43345 619321
rect 43345 619257 43409 619321
rect 43409 619257 43425 619321
rect 43425 619257 43489 619321
rect 43489 619257 43505 619321
rect 43505 619257 43516 619321
rect 42960 619177 43196 619257
rect 43280 619177 43516 619257
rect 42960 586321 43196 586413
rect 43280 586321 43516 586413
rect 42960 586257 43185 586321
rect 43185 586257 43196 586321
rect 43280 586257 43329 586321
rect 43329 586257 43345 586321
rect 43345 586257 43409 586321
rect 43409 586257 43425 586321
rect 43425 586257 43489 586321
rect 43489 586257 43505 586321
rect 43505 586257 43516 586321
rect 42960 586177 43196 586257
rect 43280 586177 43516 586257
rect 42960 553321 43196 553413
rect 43280 553321 43516 553413
rect 42960 553257 43185 553321
rect 43185 553257 43196 553321
rect 43280 553257 43329 553321
rect 43329 553257 43345 553321
rect 43345 553257 43409 553321
rect 43409 553257 43425 553321
rect 43425 553257 43489 553321
rect 43489 553257 43505 553321
rect 43505 553257 43516 553321
rect 42960 553177 43196 553257
rect 43280 553177 43516 553257
rect 42960 520321 43196 520413
rect 43280 520321 43516 520413
rect 42960 520257 43185 520321
rect 43185 520257 43196 520321
rect 43280 520257 43329 520321
rect 43329 520257 43345 520321
rect 43345 520257 43409 520321
rect 43409 520257 43425 520321
rect 43425 520257 43489 520321
rect 43489 520257 43505 520321
rect 43505 520257 43516 520321
rect 42960 520177 43196 520257
rect 43280 520177 43516 520257
rect 42960 456536 43196 456628
rect 43280 456536 43516 456628
rect 42960 456472 43185 456536
rect 43185 456472 43196 456536
rect 43280 456472 43329 456536
rect 43329 456472 43345 456536
rect 43345 456472 43409 456536
rect 43409 456472 43425 456536
rect 43425 456472 43489 456536
rect 43489 456472 43505 456536
rect 43505 456472 43516 456536
rect 42960 456392 43196 456472
rect 43280 456392 43516 456472
rect 42960 422721 43196 422813
rect 43280 422721 43516 422813
rect 42960 422657 43185 422721
rect 43185 422657 43196 422721
rect 43280 422657 43329 422721
rect 43329 422657 43345 422721
rect 43345 422657 43409 422721
rect 43409 422657 43425 422721
rect 43425 422657 43489 422721
rect 43489 422657 43505 422721
rect 43505 422657 43516 422721
rect 42960 422577 43196 422657
rect 43280 422577 43516 422657
rect 42960 389721 43196 389813
rect 43280 389721 43516 389813
rect 42960 389657 43185 389721
rect 43185 389657 43196 389721
rect 43280 389657 43329 389721
rect 43329 389657 43345 389721
rect 43345 389657 43409 389721
rect 43409 389657 43425 389721
rect 43425 389657 43489 389721
rect 43489 389657 43505 389721
rect 43505 389657 43516 389721
rect 42960 389577 43196 389657
rect 43280 389577 43516 389657
rect 42960 356464 43196 356556
rect 43280 356464 43516 356556
rect 42960 356400 43185 356464
rect 43185 356400 43196 356464
rect 43280 356400 43329 356464
rect 43329 356400 43345 356464
rect 43345 356400 43409 356464
rect 43409 356400 43425 356464
rect 43425 356400 43489 356464
rect 43489 356400 43505 356464
rect 43505 356400 43516 356464
rect 42960 356320 43196 356400
rect 43280 356320 43516 356400
rect 42960 323464 43196 323556
rect 43280 323464 43516 323556
rect 42960 323400 43185 323464
rect 43185 323400 43196 323464
rect 43280 323400 43329 323464
rect 43329 323400 43345 323464
rect 43345 323400 43409 323464
rect 43409 323400 43425 323464
rect 43425 323400 43489 323464
rect 43489 323400 43505 323464
rect 43505 323400 43516 323464
rect 42960 323320 43196 323400
rect 43280 323320 43516 323400
<< metal5 >>
rect 11127 773356 42921 773676
rect 11151 772635 43582 772676
rect 11151 772399 42960 772635
rect 43196 772399 43280 772635
rect 43516 772399 43582 772635
rect 11151 772356 43582 772399
rect 10767 771356 42921 771676
rect 10319 752366 42921 752676
rect 10448 752356 42921 752366
rect 10319 751635 43582 751676
rect 10319 751399 42960 751635
rect 43196 751399 43280 751635
rect 43516 751399 43582 751635
rect 10319 751356 43582 751399
rect 10319 750356 42921 750676
rect 9807 731356 42921 731676
rect 9807 730635 43582 730676
rect 9807 730399 42960 730635
rect 43196 730399 43280 730635
rect 43516 730399 43582 730635
rect 9807 730356 43582 730399
rect 9807 729356 42921 729676
rect 9295 710356 42921 710676
rect 9295 709635 43581 709676
rect 9295 709399 42960 709635
rect 43196 709399 43280 709635
rect 43516 709399 43581 709635
rect 9295 709356 43581 709399
rect 9295 708356 42921 708676
rect 8783 620134 42921 620454
rect 8783 619413 43581 619454
rect 8783 619177 42960 619413
rect 43196 619177 43280 619413
rect 43516 619177 43581 619413
rect 8783 619134 43581 619177
rect 8783 618134 42921 618454
rect 8271 587134 42921 587454
rect 8271 586413 43581 586454
rect 8271 586177 42960 586413
rect 43196 586177 43280 586413
rect 43516 586177 43581 586413
rect 8271 586134 43581 586177
rect 8271 585134 42921 585454
rect 7759 554134 42921 554454
rect 7759 553413 43581 553454
rect 7759 553177 42960 553413
rect 43196 553177 43280 553413
rect 43516 553177 43581 553413
rect 7759 553134 43581 553177
rect 7759 552134 42921 552454
rect 7247 521134 42921 521454
rect 7247 520413 43581 520454
rect 7247 520177 42960 520413
rect 43196 520177 43280 520413
rect 43516 520177 43581 520413
rect 7247 520134 43581 520177
rect 7247 519134 42921 519454
rect 6735 457349 42921 457669
rect 6735 456628 43581 456669
rect 6735 456392 42960 456628
rect 43196 456392 43280 456628
rect 43516 456392 43581 456628
rect 6735 456349 43581 456392
rect 6735 455349 42921 455669
rect 6223 423534 42921 423854
rect 6223 422813 43581 422854
rect 6223 422577 42960 422813
rect 43196 422577 43280 422813
rect 43516 422577 43581 422813
rect 6223 422534 43581 422577
rect 6223 421534 42921 421854
rect 5711 390534 42921 390854
rect 5711 389813 43581 389854
rect 5711 389577 42960 389813
rect 43196 389577 43280 389813
rect 43516 389577 43581 389813
rect 5711 389534 43581 389577
rect 5711 388534 42921 388854
rect 5139 357248 42921 357568
rect 42805 356568 43581 356597
rect 5139 356556 43581 356568
rect 5139 356320 42960 356556
rect 43196 356320 43280 356556
rect 43516 356320 43581 356556
rect 5139 356277 43581 356320
rect 5139 356248 43549 356277
rect 5139 355248 42921 355568
rect 4697 324277 42921 324597
rect 4697 323556 43581 323597
rect 4697 323320 42960 323556
rect 43196 323320 43280 323556
rect 43516 323320 43581 323556
rect 4697 323277 43581 323320
rect 4697 322277 42921 322597
rect 0 12000 10666 12320
rect 0 11000 10920 11320
rect 0 10000 10782 10320
rect 0 9000 10963 9320
rect 0 8000 11243 8320
rect 0 7000 11484 7320
rect 0 6000 11703 6320
rect 0 5000 12094 5320
rect 0 4000 12494 4320
rect 0 3000 12782 3320
rect 0 2000 12722 2320
rect 14521 2000 19913 2320
rect 0 1000 12858 1320
rect 14545 1000 19907 1320
rect 0 0 19133 320
use cv3_via3_30cut  cv3_via3_30cut_0
timestamp 1563083296
transform 1 0 -523607 0 1 374087
box 566656 91154 566956 91980
use cv3_via4_2cut  cv3_via4_2cut_0
timestamp 1563083296
transform 1 0 10498 0 1 772332
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_1
timestamp 1563083296
transform 1 0 9742 0 1 750324
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_2
timestamp 1563083296
transform 1 0 9245 0 1 729327
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_3
timestamp 1563083296
transform 1 0 8719 0 1 708323
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_4
timestamp 1563083296
transform 1 0 8201 0 1 618132
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_5
timestamp 1563083296
transform 1 0 7686 0 1 585114
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_6
timestamp 1563083296
transform 1 0 7173 0 1 552101
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_7
timestamp 1563083296
transform 1 0 6665 0 1 519111
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_8
timestamp 1563083296
transform 1 0 6146 0 1 455316
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_9
timestamp 1563083296
transform 1 0 5650 0 1 421519
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_10
timestamp 1563083296
transform 1 0 5148 0 1 388500
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_11
timestamp 1563083296
transform 1 0 4623 0 1 355227
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_12
timestamp 1563083296
transform 1 0 4092 0 1 322255
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_13
timestamp 1563083296
transform 1 0 13607 0 1 0
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_14
timestamp 1563083296
transform 1 0 12808 0 1 1000
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_15
timestamp 1563083296
transform 1 0 12532 0 1 1980
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_16
timestamp 1563083296
transform 1 0 12278 0 1 2986
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_17
timestamp 1563083296
transform 1 0 12020 0 1 3979
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_18
timestamp 1563083296
transform 1 0 11779 0 1 4994
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_19
timestamp 1563083296
transform 1 0 11009 0 1 7974
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_20
timestamp 1563083296
transform 1 0 19225 0 1 970
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_21
timestamp 1563083296
transform 1 0 10257 0 1 771334
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_22
timestamp 1563083296
transform 1 0 10774 0 1 773333
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_23
timestamp 1563083296
transform 1 0 9986 0 1 751348
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_24
timestamp 1563083296
transform 1 0 10240 0 1 752325
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_25
timestamp 1563083296
transform 1 0 9474 0 1 730338
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_26
timestamp 1563083296
transform 1 0 9737 0 1 731322
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_27
timestamp 1563083296
transform 1 0 8927 0 1 709332
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_28
timestamp 1563083296
transform 1 0 9229 0 1 710325
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_29
timestamp 1563083296
transform 1 0 8450 0 1 619114
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_30
timestamp 1563083296
transform 1 0 8713 0 1 620139
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_31
timestamp 1563083296
transform 1 0 7903 0 1 586113
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_32
timestamp 1563083296
transform 1 0 8223 0 1 587109
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_33
timestamp 1563083296
transform 1 0 7391 0 1 553113
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_34
timestamp 1563083296
transform 1 0 7680 0 1 554096
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_35
timestamp 1563083296
transform 1 0 6879 0 1 520113
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_36
timestamp 1563083296
transform 1 0 7179 0 1 521112
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_37
timestamp 1563083296
transform 1 0 6367 0 1 456325
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_38
timestamp 1563083296
transform 1 0 6665 0 1 457323
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_39
timestamp 1563083296
transform 1 0 5855 0 1 422513
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_40
timestamp 1563083296
transform 1 0 6146 0 1 423496
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_41
timestamp 1563083296
transform 1 0 5343 0 1 389512
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_42
timestamp 1563083296
transform 1 0 5638 0 1 390501
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_43
timestamp 1563083296
transform 1 0 4841 0 1 356224
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_44
timestamp 1563083296
transform 1 0 5113 0 1 357239
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_45
timestamp 1563083296
transform 1 0 4329 0 1 323253
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_46
timestamp 1563083296
transform 1 0 4612 0 1 324256
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_47
timestamp 1563083296
transform 1 0 13857 0 1 1000
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_48
timestamp 1563083296
transform 1 0 14133 0 1 1960
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_49
timestamp 1563083296
transform 1 0 11521 0 1 5991
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_50
timestamp 1563083296
transform 1 0 11259 0 1 6984
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_51
timestamp 1563083296
transform 1 0 10000 0 1 11983
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_52
timestamp 1563083296
transform 1 0 10742 0 1 8987
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_53
timestamp 1563083296
transform 1 0 10496 0 1 9978
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_54
timestamp 1563083296
transform 1 0 10250 0 1 10974
box 0 0 688 368
<< properties >>
string FIXED_BBOX 0 0 44160 800234
<< end >>
