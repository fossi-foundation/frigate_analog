magic
tech sky130A
magscale 1 2
timestamp 1719932489
<< isosubstrate >>
rect 284 560 3656 3458
<< viali >>
rect 1663 2610 1697 2644
rect 1951 2610 1985 2644
rect 2431 1944 2465 1978
<< metal1 >>
rect 480 3282 3456 3307
rect 480 3230 2122 3282
rect 2174 3230 2186 3282
rect 2238 3230 3456 3282
rect 480 3205 3456 3230
rect 1651 2644 1709 2650
rect 1651 2610 1663 2644
rect 1697 2641 1709 2644
rect 1939 2644 1997 2650
rect 1939 2641 1951 2644
rect 1697 2613 1951 2641
rect 1697 2610 1709 2613
rect 1651 2604 1709 2610
rect 1939 2610 1951 2613
rect 1985 2641 1997 2644
rect 3184 2641 3190 2653
rect 1985 2613 3190 2641
rect 1985 2610 1997 2613
rect 1939 2604 1997 2610
rect 3184 2601 3190 2613
rect 3242 2601 3248 2653
rect 480 2468 3456 2493
rect 480 2416 822 2468
rect 874 2416 886 2468
rect 938 2416 3456 2468
rect 480 2391 3456 2416
rect 1536 2286 2110 2289
rect 1536 2232 1670 2286
rect 1664 2226 1670 2232
rect 1854 2232 2110 2286
rect 1854 2226 1860 2232
rect 1664 2222 1860 2226
rect 592 1935 598 1987
rect 650 1975 656 1987
rect 2419 1978 2477 1984
rect 2419 1975 2431 1978
rect 650 1947 2431 1975
rect 650 1935 656 1947
rect 2419 1944 2431 1947
rect 2465 1944 2477 1978
rect 2419 1938 2477 1944
rect 480 1654 3456 1679
rect 480 1602 2122 1654
rect 2174 1602 2186 1654
rect 2238 1602 3456 1654
rect 480 1577 3456 1602
rect 480 840 3456 865
rect 480 788 822 840
rect 874 788 886 840
rect 938 788 3456 840
rect 480 763 3456 788
<< via1 >>
rect 2122 3230 2174 3282
rect 2186 3230 2238 3282
rect 3190 2601 3242 2653
rect 822 2416 874 2468
rect 886 2416 938 2468
rect 1670 2226 1854 2286
rect 598 1935 650 1987
rect 2122 1602 2174 1654
rect 2186 1602 2238 1654
rect 822 788 874 840
rect 886 788 938 840
<< metal2 >>
rect 2112 3284 2248 3307
rect 2168 3282 2192 3284
rect 2174 3230 2186 3282
rect 2168 3228 2192 3230
rect 2112 3205 2248 3228
rect 3190 2653 3242 2659
rect 3284 2604 3340 3800
rect 3242 2601 3340 2604
rect 3190 2600 3340 2601
rect 3190 2595 3326 2600
rect 3202 2576 3326 2595
rect 812 2470 948 2493
rect 868 2468 892 2470
rect 874 2416 886 2468
rect 868 2414 892 2416
rect 812 2391 948 2414
rect 1660 2286 1864 2296
rect 1660 2226 1670 2286
rect 1854 2226 1864 2286
rect 1660 2214 1864 2226
rect 598 1987 650 1993
rect 598 1929 650 1935
rect 610 800 638 1929
rect 2112 1656 2248 1679
rect 2168 1654 2192 1656
rect 2174 1602 2186 1654
rect 2168 1600 2192 1602
rect 2112 1577 2248 1600
rect 812 842 948 865
rect 868 840 892 842
rect 596 -400 652 800
rect 874 788 886 840
rect 868 786 892 788
rect 812 763 948 786
<< via2 >>
rect 2112 3282 2168 3284
rect 2192 3282 2248 3284
rect 2112 3230 2122 3282
rect 2122 3230 2168 3282
rect 2192 3230 2238 3282
rect 2238 3230 2248 3282
rect 2112 3228 2168 3230
rect 2192 3228 2248 3230
rect 812 2468 868 2470
rect 892 2468 948 2470
rect 812 2416 822 2468
rect 822 2416 868 2468
rect 892 2416 938 2468
rect 938 2416 948 2468
rect 812 2414 868 2416
rect 892 2414 948 2416
rect 1670 2226 1854 2286
rect 2112 1654 2168 1656
rect 2192 1654 2248 1656
rect 2112 1602 2122 1654
rect 2122 1602 2168 1654
rect 2192 1602 2238 1654
rect 2238 1602 2248 1654
rect 2112 1600 2168 1602
rect 2192 1600 2248 1602
rect 812 840 868 842
rect 892 840 948 842
rect 812 788 822 840
rect 822 788 868 840
rect 892 788 938 840
rect 938 788 948 840
rect 812 786 868 788
rect 892 786 948 788
<< metal3 >>
rect 2090 3288 2270 3289
rect 2090 3224 2108 3288
rect 2172 3224 2188 3288
rect 2252 3224 2270 3288
rect 2090 3223 2270 3224
rect 790 2474 970 2475
rect 790 2410 808 2474
rect 872 2410 888 2474
rect 952 2410 970 2474
rect 790 2409 970 2410
rect 1660 2290 1864 2296
rect 1660 2226 1670 2290
rect 1854 2226 1864 2290
rect 1660 2214 1864 2226
rect 2090 1660 2270 1661
rect 2090 1596 2108 1660
rect 2172 1596 2188 1660
rect 2252 1596 2270 1660
rect 2090 1595 2270 1596
rect 790 846 970 847
rect 790 782 808 846
rect 872 782 888 846
rect 952 782 970 846
rect 790 781 970 782
<< via3 >>
rect 2108 3284 2172 3288
rect 2108 3228 2112 3284
rect 2112 3228 2168 3284
rect 2168 3228 2172 3284
rect 2108 3224 2172 3228
rect 2188 3284 2252 3288
rect 2188 3228 2192 3284
rect 2192 3228 2248 3284
rect 2248 3228 2252 3284
rect 2188 3224 2252 3228
rect 808 2470 872 2474
rect 808 2414 812 2470
rect 812 2414 868 2470
rect 868 2414 872 2470
rect 808 2410 872 2414
rect 888 2470 952 2474
rect 888 2414 892 2470
rect 892 2414 948 2470
rect 948 2414 952 2470
rect 888 2410 952 2414
rect 1670 2286 1854 2290
rect 1670 2226 1854 2286
rect 2108 1656 2172 1660
rect 2108 1600 2112 1656
rect 2112 1600 2168 1656
rect 2168 1600 2172 1656
rect 2108 1596 2172 1600
rect 2188 1656 2252 1660
rect 2188 1600 2192 1656
rect 2192 1600 2248 1656
rect 2248 1600 2252 1656
rect 2188 1596 2252 1600
rect 808 842 872 846
rect 808 786 812 842
rect 812 786 868 842
rect 868 786 872 842
rect 808 782 872 786
rect 888 842 952 846
rect 888 786 892 842
rect 892 786 948 842
rect 948 786 952 842
rect 888 782 952 786
<< metal4 >>
rect 790 2474 970 3307
rect 2090 3288 2270 3307
rect 790 2410 808 2474
rect 872 2410 888 2474
rect 952 2410 970 2474
rect 790 846 970 2410
rect 1670 2296 1850 3256
rect 2090 3224 2108 3288
rect 2172 3224 2188 3288
rect 2252 3224 2270 3288
rect 1660 2290 1860 2296
rect 1660 2226 1670 2290
rect 1854 2226 1860 2290
rect 1660 2216 1860 2226
rect 790 782 808 846
rect 872 782 888 846
rect 952 782 970 846
rect 1670 814 1850 2216
rect 2090 1660 2270 3224
rect 2090 1596 2108 1660
rect 2172 1596 2188 1660
rect 2252 1596 2270 1660
rect 790 763 970 782
rect 2090 763 2270 1596
rect 2970 814 3150 3256
use sky130_fd_sc_hvl__diode_2  ANTENNA_lvlshiftdown_A $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 1536 0 -1 3256
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 480 0 -1 1628
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_8
timestamp 1715205430
transform 1 0 1248 0 -1 1628
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_16
timestamp 1715205430
transform 1 0 2016 0 -1 1628
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 2784 0 -1 1628
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_0_28 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 3168 0 -1 1628
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_1  FILLER_0_30 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 3360 0 -1 1628
box -66 -43 162 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_0
timestamp 1715205430
transform 1 0 480 0 1 1628
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_1_8
timestamp 1715205430
transform 1 0 1248 0 1 1628
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_1  FILLER_1_12
timestamp 1715205430
transform 1 0 1632 0 1 1628
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  FILLER_1_30
timestamp 1715205430
transform 1 0 3360 0 1 1628
box -66 -43 162 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_0
timestamp 1715205430
transform 1 0 480 0 -1 3256
box -66 -43 834 897
use sky130_fd_sc_hvl__fill_2  FILLER_2_8
timestamp 1715205430
transform 1 0 1248 0 -1 3256
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_1  FILLER_2_10
timestamp 1715205430
transform 1 0 1440 0 -1 3256
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  FILLER_2_30
timestamp 1715205430
transform 1 0 3360 0 -1 3256
box -66 -43 162 897
use sky130_fd_sc_hvl__lsbufhv2lv_1  lvlshiftdown $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1715205430
transform 1 0 1728 0 1 1628
box -66 -43 1698 1671
<< labels >>
rlabel metal2 s 3284 2600 3340 3800 6 A
port 0 nsew signal input
rlabel metal2 s 596 -400 652 800 6 X
port 1 nsew signal tristate
rlabel metal4 s 790 763 970 3307 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 2090 763 2270 3307 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 1670 814 1850 3256 6 LVPWR
port 4 nsew power bidirectional
rlabel metal4 s 2970 814 3150 3256 6 LVGND
port 5 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 4000 3400
<< end >>
