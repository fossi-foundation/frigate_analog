magic
tech sky130A
magscale 1 2
timestamp 1717859897
<< metal2 >>
rect 630 31091 944 31117
rect 630 30712 663 31091
rect 912 30712 944 31091
rect 630 30683 944 30712
<< via2 >>
rect 663 30712 912 31091
<< metal3 >>
rect 600 31092 1050 31117
rect 600 30676 628 31092
rect 1022 30676 1050 31092
rect 600 30642 1050 30676
<< via3 >>
rect 628 31091 1022 31092
rect 628 30712 663 31091
rect 663 30712 912 31091
rect 912 30712 1022 31091
rect 628 30676 1022 30712
<< metal4 >>
rect 600 31092 1050 31117
rect 600 30676 628 31092
rect 1022 30676 1050 31092
rect 600 30642 1050 30676
rect 0 949 200 30415
rect 0 905 320 949
rect 0 194 38 905
rect 279 194 320 905
rect 0 149 320 194
rect 600 0 800 30642
rect 1200 949 1400 30420
rect 1080 903 1400 949
rect 1080 192 1121 903
rect 1362 192 1400 903
rect 1080 149 1400 192
<< via4 >>
rect 38 194 279 905
rect 1121 192 1362 903
<< metal5 >>
rect 0 905 1401 949
rect 0 194 38 905
rect 279 903 1401 905
rect 279 194 1121 903
rect 0 192 1121 194
rect 1362 192 1401 903
rect 0 149 1401 192
<< properties >>
string FIXED_BBOX 0 0 1401 31117
string LEFclass COVER
<< end >>
