magic
tech sky130A
magscale 1 2
timestamp 1721093827
<< metal4 >>
rect -1349 1039 1349 1080
rect -1349 -1039 1093 1039
rect 1329 -1039 1349 1039
rect -1349 -1080 1349 -1039
<< via4 >>
rect 1093 -1039 1329 1039
<< mimcap2 >>
rect -1269 960 731 1000
rect -1269 -960 -1229 960
rect 691 -960 731 960
rect -1269 -1000 731 -960
<< mimcap2contact >>
rect -1229 -960 691 960
<< metal5 >>
rect 1051 1039 1371 1081
rect -1253 960 715 984
rect -1253 -960 -1229 960
rect 691 -960 715 960
rect -1253 -984 715 -960
rect 1051 -1039 1093 1039
rect 1329 -1039 1371 1039
rect 1051 -1081 1371 -1039
<< properties >>
string FIXED_BBOX -1349 -1080 811 1080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 10.00 l 10.00 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
