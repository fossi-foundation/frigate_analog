magic
tech sky130A
magscale 1 2
timestamp 1719433677
<< checkpaint >>
rect 431918 70502 432946 70630
<< metal3 >>
rect 431918 70623 432946 70630
rect 431918 70510 431928 70623
rect 432938 70510 432946 70623
rect 431918 70502 432946 70510
<< via3 >>
rect 431928 70510 432938 70623
<< metal4 >>
rect 431918 70623 432946 70630
rect 431918 70510 431928 70623
rect 432938 70510 432946 70623
rect 431918 70502 432946 70510
<< end >>
