magic
tech sky130A
magscale 1 2
timestamp 1724444338
<< metal1 >>
rect -214 2415 -208 2467
rect -156 2459 -150 2467
rect -156 2423 30 2459
rect -156 2415 -150 2423
rect 4302 2415 4308 2467
rect 4360 2459 4366 2467
rect 4360 2423 4546 2459
rect 4360 2415 4366 2423
rect 8818 2415 8824 2467
rect 8876 2459 8882 2467
rect 8876 2423 9062 2459
rect 8876 2415 8882 2423
rect 15788 2411 15794 2463
rect 15846 2455 15852 2463
rect 15846 2419 16010 2455
rect 15846 2411 15852 2419
rect 20304 2411 20310 2463
rect 20362 2455 20368 2463
rect 20362 2419 20526 2455
rect 20362 2411 20368 2419
rect 24820 2411 24826 2463
rect 24878 2455 24884 2463
rect 24878 2419 25040 2455
rect 24878 2411 24884 2419
rect 4 2007 298 2018
rect 4 1891 18 2007
rect 276 1891 298 2007
rect 4520 2007 4814 2018
rect 4520 1891 4534 2007
rect 4792 1891 4814 2007
rect 9036 2007 9330 2018
rect 9036 1891 9050 2007
rect 9308 1891 9330 2007
rect 16046 2014 16340 2025
rect 16046 1897 16060 2014
rect 16318 1897 16340 2014
rect 16046 1891 16340 1897
rect 20562 2014 20856 2025
rect 20562 1897 20576 2014
rect 20834 1897 20856 2014
rect 20562 1891 20856 1897
rect 25078 2014 25372 2025
rect 25078 1897 25092 2014
rect 25350 1897 25372 2014
rect 25078 1891 25372 1897
<< via1 >>
rect 2536 2492 3050 2561
rect 7052 2492 7566 2561
rect 11568 2492 12082 2561
rect 18578 2499 19092 2568
rect 23094 2499 23608 2568
rect 27610 2499 28124 2568
rect -208 2415 -156 2467
rect 4308 2415 4360 2467
rect 8824 2415 8876 2467
rect 15794 2411 15846 2463
rect 20310 2411 20362 2463
rect 24826 2411 24878 2463
rect 18 1891 276 2007
rect 4534 1891 4792 2007
rect 9050 1891 9308 2007
rect 16060 1897 16318 2014
rect 20576 1897 20834 2014
rect 25092 1897 25350 2014
<< metal2 >>
rect 406 4121 13503 4551
rect -664 3555 414 3991
rect 3852 3555 4930 3991
rect 8368 3555 9446 3991
rect -664 869 -308 3555
rect 2517 2566 3065 2579
rect 2517 2561 2537 2566
rect 2517 2492 2536 2561
rect -208 2467 -156 2473
rect 2517 2460 2537 2492
rect 3054 2460 3065 2566
rect 2517 2448 3065 2460
rect -208 2409 -156 2415
rect -200 883 -164 2409
rect 4 2007 298 2018
rect 4 1890 18 2007
rect 276 1890 298 2007
rect 4 1877 298 1890
rect 3852 869 4208 3555
rect 7033 2566 7581 2579
rect 7033 2561 7053 2566
rect 7033 2492 7052 2561
rect 4308 2467 4360 2473
rect 7033 2460 7053 2492
rect 7570 2460 7581 2566
rect 7033 2448 7581 2460
rect 4308 2409 4360 2415
rect 4316 883 4352 2409
rect 4520 2007 4814 2018
rect 4520 1890 4534 2007
rect 4792 1890 4814 2007
rect 4520 1877 4814 1890
rect 8368 869 8724 3555
rect 11549 2566 12097 2579
rect 11549 2561 11569 2566
rect 11549 2492 11568 2561
rect 8824 2467 8876 2473
rect 11549 2460 11569 2492
rect 12086 2460 12097 2566
rect 11549 2448 12097 2460
rect 8824 2409 8876 2415
rect 8832 883 8868 2409
rect 9036 2007 9330 2018
rect 9036 1890 9050 2007
rect 9308 1890 9330 2007
rect 9036 1877 9330 1890
rect 13073 858 13503 4121
rect 15127 4123 28524 4553
rect 15127 858 15557 4123
rect 19482 3559 20156 3989
rect 18559 2573 19107 2586
rect 18559 2568 18579 2573
rect 18559 2499 18578 2568
rect 15794 2463 15846 2469
rect 18559 2467 18579 2499
rect 19096 2467 19107 2573
rect 18559 2455 19107 2467
rect 15794 2405 15846 2411
rect 15802 887 15838 2405
rect 16046 2014 16340 2025
rect 16046 1897 16060 2014
rect 16318 1897 16340 2014
rect 16046 1884 16340 1897
rect 19800 867 20156 3559
rect 23984 3559 24672 3989
rect 23984 3557 24010 3559
rect 23075 2573 23623 2586
rect 23075 2568 23095 2573
rect 23075 2499 23094 2568
rect 20310 2463 20362 2469
rect 23075 2467 23095 2499
rect 23612 2467 23623 2573
rect 23075 2455 23623 2467
rect 20310 2405 20362 2411
rect 20318 887 20354 2405
rect 20562 2014 20856 2025
rect 20562 1897 20576 2014
rect 20834 1897 20856 2014
rect 20562 1884 20856 1897
rect 24316 867 24672 3559
rect 28500 3559 29188 3989
rect 28500 3557 28526 3559
rect 27591 2573 28139 2586
rect 27591 2568 27611 2573
rect 27591 2499 27610 2568
rect 24826 2463 24878 2469
rect 27591 2467 27611 2499
rect 28128 2467 28139 2573
rect 27591 2455 28139 2467
rect 24826 2405 24878 2411
rect 24834 887 24870 2405
rect 25078 2014 25372 2025
rect 25078 1897 25092 2014
rect 25350 1897 25372 2014
rect 25078 1884 25372 1897
rect 28832 867 29188 3559
<< via2 >>
rect 640 4718 1542 4854
rect 5156 4718 6058 4854
rect 9672 4718 10574 4854
rect 16682 4725 17584 4861
rect 21198 4725 22100 4861
rect 25714 4725 26616 4861
rect 673 3253 1575 3389
rect 2537 2561 3054 2566
rect 2537 2492 3050 2561
rect 3050 2492 3054 2561
rect 2537 2460 3054 2492
rect 18 1891 276 2007
rect 18 1890 276 1891
rect 5189 3253 6091 3389
rect 7053 2561 7570 2566
rect 7053 2492 7566 2561
rect 7566 2492 7570 2561
rect 7053 2460 7570 2492
rect 4534 1891 4792 2007
rect 4534 1890 4792 1891
rect 9705 3253 10607 3389
rect 11569 2561 12086 2566
rect 11569 2492 12082 2561
rect 12082 2492 12086 2561
rect 11569 2460 12086 2492
rect 9050 1891 9308 2007
rect 9050 1890 9308 1891
rect 16715 3260 17617 3396
rect 18579 2568 19096 2573
rect 18579 2499 19092 2568
rect 19092 2499 19096 2568
rect 18579 2467 19096 2499
rect 16060 1897 16318 2014
rect 21231 3260 22133 3396
rect 23095 2568 23612 2573
rect 23095 2499 23608 2568
rect 23608 2499 23612 2568
rect 23095 2467 23612 2499
rect 20576 1897 20834 2014
rect 25747 3260 26649 3396
rect 27611 2568 28128 2573
rect 27611 2499 28124 2568
rect 28124 2499 28128 2568
rect 27611 2467 28128 2499
rect 25092 1897 25350 2014
<< metal3 >>
rect 16588 4869 17683 4876
rect 21104 4869 22199 4876
rect 25620 4869 26715 4876
rect -14 4861 28516 4869
rect -14 4854 16682 4861
rect -14 4718 640 4854
rect 1542 4718 5156 4854
rect 6058 4718 9672 4854
rect 10574 4725 16682 4854
rect 17584 4725 21198 4861
rect 22100 4725 25714 4861
rect 26616 4725 28516 4861
rect 10574 4718 28516 4725
rect -14 4700 28516 4718
rect 16616 3405 17711 3412
rect 21132 3405 22227 3412
rect 25648 3405 26743 3412
rect -14 3396 28516 3405
rect -14 3389 16715 3396
rect -14 3253 673 3389
rect 1575 3253 5189 3389
rect 6091 3253 9705 3389
rect 10607 3260 16715 3389
rect 17617 3260 21231 3396
rect 22133 3260 25747 3396
rect 26649 3260 28516 3396
rect 10607 3253 28516 3260
rect -14 3236 28516 3253
rect 18446 2599 19271 2606
rect 22962 2599 23787 2606
rect 27478 2599 28303 2606
rect 47 2573 28577 2599
rect 47 2566 18579 2573
rect 47 2460 2537 2566
rect 3054 2460 7053 2566
rect 7570 2460 11569 2566
rect 12086 2467 18579 2566
rect 19096 2467 23095 2573
rect 23612 2467 27611 2573
rect 28128 2467 28577 2573
rect 12086 2460 28577 2467
rect 47 2430 28577 2460
rect 16035 2030 16440 2037
rect 20551 2030 20956 2037
rect 25067 2030 25472 2037
rect -7 2014 28523 2030
rect -7 2007 16060 2014
rect -7 1890 18 2007
rect 276 1890 4534 2007
rect 4792 1890 9050 2007
rect 9308 1897 16060 2007
rect 16318 1897 20576 2014
rect 20834 1897 25092 2014
rect 25350 1897 28523 2014
rect 9308 1890 28523 1897
rect -7 1861 28523 1890
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_0 ../ip/sky130_ef_ip__analog_switches/mag
array 0 2 4516 0 0 -4248
timestamp 1724439637
transform 1 0 0 0 -1 4529
box -4 -600 3538 3648
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_1
array 0 2 4516 0 0 -4248
timestamp 1724439637
transform 1 0 16000 0 -1 4529
box -4 -600 3538 3648
<< end >>
