magic
tech sky130A
timestamp 1719247715
<< checkpaint >>
rect 7167 52462 7297 52805
<< metal1 >>
rect 7167 52791 7297 52805
rect 7167 52475 7181 52791
rect 7286 52475 7297 52791
rect 7167 52462 7297 52475
<< via1 >>
rect 7181 52475 7286 52791
<< metal2 >>
rect 7167 52791 7297 52805
rect 7167 52475 7181 52791
rect 7286 52475 7297 52791
rect 7167 52462 7297 52475
<< end >>
