VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_routes_top
  CLASS COVER ;
  FOREIGN analog_routes_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.000 BY 154.845 ;
  OBS
      LAYER met2 ;
        RECT 0.655 153.150 2.465 154.845 ;
        RECT 3.745 153.150 7.000 154.845 ;
      LAYER met3 ;
        RECT 0.655 153.150 3.000 154.845 ;
        RECT 4.655 153.150 7.000 154.845 ;
      LAYER met4 ;
        RECT 0.655 153.150 3.000 154.845 ;
        RECT 4.655 153.150 7.000 154.845 ;
        RECT 0.000 0.000 1.000 152.230 ;
        RECT 2.000 0.000 3.000 153.150 ;
        RECT 4.000 0.000 5.000 152.230 ;
        RECT 6.000 0.000 7.000 153.150 ;
        RECT 8.000 0.000 9.000 152.230 ;
  END
END analog_routes_top
END LIBRARY

