magic
tech sky130A
magscale 1 2
timestamp 1719257891
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_1 ../dependencies/sky130_ef_ip__analog_switches/mag
array 0 2 -4515 0 3 -4632
timestamp 1719257891
transform 0 -1 3580 -1 0 4419
box -4 -600 3538 3648
<< end >>
