VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_routes_right
  CLASS COVER ;
  FOREIGN analog_routes_right ;
  ORIGIN 0.000 0.000 ;
  SIZE 220.800 BY 4001.170 ;
  OBS
      LAYER met2 ;
        RECT 221.840 2933.575 222.080 2944.825 ;
        RECT 221.840 2768.485 222.080 2779.685 ;
        RECT 221.840 2603.505 222.080 2614.745 ;
        RECT 221.840 2440.175 222.080 2449.875 ;
        RECT 220.695 2439.935 222.080 2440.175 ;
        RECT 217.205 2329.235 218.475 2329.665 ;
        RECT 220.695 2329.235 220.935 2439.935 ;
        RECT 217.205 2328.995 220.935 2329.235 ;
        RECT 217.205 2328.415 218.475 2328.995 ;
        RECT 214.895 2282.415 220.995 2282.655 ;
        RECT 214.895 2138.095 215.135 2282.415 ;
        RECT 214.895 2137.855 222.080 2138.095 ;
        RECT 221.840 2115.635 222.080 2137.855 ;
        RECT 221.840 1950.635 222.080 1961.825 ;
        RECT 221.840 1785.455 222.080 1796.805 ;
        RECT 221.840 1620.665 222.080 1631.705 ;
        RECT 98.195 1.930 99.535 4.705 ;
      LAYER met3 ;
        RECT 215.760 3862.230 219.590 3862.875 ;
        RECT 215.760 3757.230 219.590 3757.875 ;
        RECT 215.760 3652.230 219.590 3652.875 ;
        RECT 215.760 3547.230 219.590 3547.875 ;
        RECT 215.760 3096.720 219.590 3096.765 ;
        RECT 215.760 3096.120 220.800 3096.720 ;
        RECT 215.760 2931.720 219.590 2931.765 ;
        RECT 215.760 2931.120 220.800 2931.720 ;
        RECT 215.760 2766.720 219.590 2766.765 ;
        RECT 215.760 2766.120 220.800 2766.720 ;
        RECT 215.760 2601.720 219.590 2601.765 ;
        RECT 215.760 2601.120 220.800 2601.720 ;
        RECT 215.245 2330.120 216.745 2330.335 ;
        RECT 215.245 2328.120 219.475 2330.120 ;
        RECT 215.245 2326.205 216.745 2328.120 ;
        RECT 215.760 2282.795 219.590 2282.840 ;
        RECT 215.760 2282.195 220.800 2282.795 ;
        RECT 215.760 2113.720 219.590 2113.765 ;
        RECT 215.760 2113.120 220.800 2113.720 ;
        RECT 215.760 1948.720 219.590 1948.765 ;
        RECT 215.760 1948.120 220.800 1948.720 ;
        RECT 215.760 1782.435 219.590 1782.480 ;
        RECT 215.760 1781.835 220.800 1782.435 ;
        RECT 215.760 1617.435 219.590 1617.480 ;
        RECT 215.760 1616.835 220.800 1617.435 ;
        RECT 97.655 1.930 99.530 5.000 ;
      LAYER met4 ;
        RECT 2.675 1587.405 3.315 4001.170 ;
        RECT 3.975 1588.705 4.615 4001.170 ;
        RECT 5.235 1589.965 5.875 4001.170 ;
        RECT 6.535 1591.265 7.175 4001.170 ;
        RECT 7.795 1592.525 8.435 4001.170 ;
        RECT 9.095 1593.825 9.735 4001.170 ;
        RECT 10.355 1595.085 10.995 4001.170 ;
        RECT 11.655 1596.385 12.295 4001.170 ;
        RECT 12.915 1597.645 13.555 4001.170 ;
        RECT 14.215 1598.945 14.855 4001.170 ;
        RECT 15.475 1600.205 16.115 4001.170 ;
        RECT 16.775 1601.505 17.415 4001.170 ;
        RECT 18.035 1602.765 18.675 4001.170 ;
        RECT 19.335 1604.065 19.975 4001.170 ;
        RECT 20.595 1612.995 21.235 4001.170 ;
        RECT 21.895 1617.985 22.535 4001.170 ;
        RECT 23.195 1777.855 23.835 4001.170 ;
        RECT 24.455 1782.840 25.095 4001.170 ;
        RECT 25.755 1944.220 26.395 4001.170 ;
        RECT 27.015 1949.280 27.655 4001.170 ;
        RECT 28.315 2109.315 28.955 4001.170 ;
        RECT 29.575 2114.285 30.215 4001.170 ;
        RECT 30.875 2278.300 31.515 4001.170 ;
        RECT 32.135 2283.345 32.775 4001.170 ;
        RECT 33.435 2597.275 34.075 4001.170 ;
        RECT 34.695 2602.285 35.335 4001.170 ;
        RECT 35.995 2762.225 36.635 4001.170 ;
        RECT 37.255 2767.285 37.895 4001.170 ;
        RECT 38.555 2927.290 39.195 4001.170 ;
        RECT 39.815 2932.285 40.455 4001.170 ;
        RECT 41.115 3092.380 41.755 4001.170 ;
        RECT 42.375 3097.290 43.015 4001.170 ;
        RECT 43.675 3543.335 44.315 4001.170 ;
        RECT 44.935 3548.380 45.575 4001.170 ;
        RECT 46.235 3648.355 46.875 4001.170 ;
        RECT 47.495 3653.410 48.135 4001.170 ;
        RECT 48.795 3753.340 49.435 4001.170 ;
        RECT 50.055 3758.460 50.695 4001.170 ;
        RECT 51.355 3858.390 51.995 4001.170 ;
        RECT 52.615 3863.380 53.255 4001.170 ;
        RECT 53.915 3868.385 54.555 4001.170 ;
        RECT 53.915 3867.125 57.190 3868.385 ;
        RECT 53.990 3866.785 57.190 3867.125 ;
        RECT 52.610 3861.780 55.810 3863.380 ;
        RECT 214.460 3862.875 217.905 3863.380 ;
        RECT 214.460 3862.230 219.590 3862.875 ;
        RECT 214.460 3861.780 217.905 3862.230 ;
        RECT 51.355 3856.790 54.605 3858.390 ;
        RECT 51.355 3763.345 51.995 3856.790 ;
        RECT 51.320 3761.745 54.520 3763.345 ;
        RECT 50.050 3756.860 53.250 3758.460 ;
        RECT 214.460 3757.875 217.905 3758.380 ;
        RECT 214.460 3757.230 219.590 3757.875 ;
        RECT 214.460 3756.780 217.905 3757.230 ;
        RECT 48.795 3751.740 52.030 3753.340 ;
        RECT 48.795 3658.330 49.435 3751.740 ;
        RECT 48.795 3656.730 52.005 3658.330 ;
        RECT 48.795 3656.485 49.435 3656.730 ;
        RECT 47.490 3651.810 50.690 3653.410 ;
        RECT 214.460 3652.875 217.905 3653.380 ;
        RECT 214.460 3652.230 219.590 3652.875 ;
        RECT 214.460 3651.780 217.905 3652.230 ;
        RECT 46.235 3646.755 49.545 3648.355 ;
        RECT 46.235 3553.345 46.875 3646.755 ;
        RECT 46.235 3551.745 49.465 3553.345 ;
        RECT 46.235 3551.595 46.875 3551.745 ;
        RECT 44.755 3546.780 47.955 3548.380 ;
        RECT 214.460 3547.875 217.905 3548.380 ;
        RECT 214.460 3547.230 219.590 3547.875 ;
        RECT 214.460 3546.780 217.905 3547.230 ;
        RECT 43.675 3541.735 46.915 3543.335 ;
        RECT 43.675 3102.415 44.315 3541.735 ;
        RECT 43.675 3100.815 46.885 3102.415 ;
        RECT 43.675 3100.730 44.315 3100.815 ;
        RECT 42.370 3095.690 45.570 3097.290 ;
        RECT 214.460 3096.765 217.905 3097.270 ;
        RECT 214.460 3096.120 219.590 3096.765 ;
        RECT 214.460 3095.670 217.905 3096.120 ;
        RECT 41.115 3090.780 44.325 3092.380 ;
        RECT 41.115 2937.265 41.755 3090.780 ;
        RECT 41.115 2935.665 44.435 2937.265 ;
        RECT 41.115 2935.415 41.755 2935.665 ;
        RECT 39.635 2930.685 42.835 2932.285 ;
        RECT 214.460 2931.765 217.905 2932.270 ;
        RECT 214.460 2931.120 219.590 2931.765 ;
        RECT 214.460 2930.670 217.905 2931.120 ;
        RECT 38.550 2925.690 41.750 2927.290 ;
        RECT 38.555 2772.200 39.195 2925.690 ;
        RECT 38.520 2770.600 41.720 2772.200 ;
        RECT 37.075 2765.685 40.275 2767.285 ;
        RECT 214.460 2766.765 217.905 2767.270 ;
        RECT 214.460 2766.120 219.590 2766.765 ;
        RECT 214.460 2765.670 217.905 2766.120 ;
        RECT 35.985 2760.625 39.185 2762.225 ;
        RECT 35.995 2607.280 36.635 2760.625 ;
        RECT 35.995 2605.680 39.215 2607.280 ;
        RECT 35.995 2605.120 36.635 2605.680 ;
        RECT 34.515 2600.685 37.715 2602.285 ;
        RECT 214.460 2601.765 217.905 2602.270 ;
        RECT 214.460 2601.120 219.590 2601.765 ;
        RECT 214.460 2600.670 217.905 2601.120 ;
        RECT 33.435 2595.675 36.645 2597.275 ;
        RECT 33.435 2288.335 34.075 2595.675 ;
        RECT 215.645 2330.335 216.405 2330.365 ;
        RECT 215.245 2326.205 216.745 2330.335 ;
        RECT 33.435 2286.735 36.645 2288.335 ;
        RECT 33.435 2286.120 34.075 2286.735 ;
        RECT 215.645 2283.345 216.405 2326.205 ;
        RECT 31.955 2281.745 35.155 2283.345 ;
        RECT 214.460 2282.840 217.905 2283.345 ;
        RECT 214.460 2282.195 219.590 2282.840 ;
        RECT 214.460 2281.745 217.905 2282.195 ;
        RECT 30.850 2276.700 34.050 2278.300 ;
        RECT 30.875 2119.200 31.515 2276.700 ;
        RECT 30.850 2117.600 34.050 2119.200 ;
        RECT 30.875 2117.245 31.515 2117.600 ;
        RECT 29.395 2112.685 32.595 2114.285 ;
        RECT 214.460 2113.765 217.905 2114.270 ;
        RECT 214.460 2113.120 219.590 2113.765 ;
        RECT 214.460 2112.670 217.905 2113.120 ;
        RECT 28.315 2107.715 31.570 2109.315 ;
        RECT 28.315 1954.225 28.955 2107.715 ;
        RECT 28.310 1952.625 31.510 1954.225 ;
        RECT 28.315 1952.435 28.955 1952.625 ;
        RECT 26.835 1947.680 30.035 1949.280 ;
        RECT 214.460 1948.765 217.905 1949.270 ;
        RECT 214.460 1948.120 219.590 1948.765 ;
        RECT 214.460 1947.670 217.905 1948.120 ;
        RECT 25.755 1942.620 29.060 1944.220 ;
        RECT 25.755 1787.915 26.395 1942.620 ;
        RECT 25.685 1786.315 28.885 1787.915 ;
        RECT 24.325 1781.240 27.525 1782.840 ;
        RECT 214.460 1782.480 217.905 1782.985 ;
        RECT 214.460 1781.835 219.590 1782.480 ;
        RECT 214.460 1781.385 217.905 1781.835 ;
        RECT 23.195 1776.255 26.435 1777.855 ;
        RECT 23.195 1623.000 23.835 1776.255 ;
        RECT 23.180 1621.400 26.380 1623.000 ;
        RECT 21.765 1616.385 24.965 1617.985 ;
        RECT 214.460 1617.480 217.905 1617.985 ;
        RECT 214.460 1616.835 219.590 1617.480 ;
        RECT 214.460 1616.385 217.905 1616.835 ;
        RECT 20.580 1611.395 23.780 1612.995 ;
        RECT 20.595 1605.325 21.235 1611.395 ;
        RECT 20.595 1604.685 71.235 1605.325 ;
        RECT 19.335 1603.425 69.975 1604.065 ;
        RECT 18.035 1602.125 68.675 1602.765 ;
        RECT 16.775 1600.865 67.415 1601.505 ;
        RECT 15.475 1599.565 66.115 1600.205 ;
        RECT 14.215 1598.305 64.855 1598.945 ;
        RECT 12.915 1597.005 63.555 1597.645 ;
        RECT 11.655 1595.745 62.295 1596.385 ;
        RECT 10.355 1594.445 60.995 1595.085 ;
        RECT 9.095 1593.185 59.735 1593.825 ;
        RECT 7.795 1591.885 58.435 1592.525 ;
        RECT 6.535 1590.625 57.175 1591.265 ;
        RECT 5.235 1589.325 55.875 1589.965 ;
        RECT 3.975 1588.065 54.615 1588.705 ;
        RECT 52.675 1587.405 53.315 1587.410 ;
        RECT 2.675 1586.780 53.315 1587.405 ;
        RECT 31.370 1586.765 53.315 1586.780 ;
        RECT 52.675 61.635 53.315 1586.765 ;
        RECT 50.120 60.035 53.320 61.635 ;
        RECT 53.975 56.590 54.615 1588.065 ;
        RECT 51.370 55.900 54.615 56.590 ;
        RECT 51.370 54.990 54.570 55.900 ;
        RECT 55.235 51.610 55.875 1589.325 ;
        RECT 52.600 50.615 55.875 51.610 ;
        RECT 52.600 50.010 55.800 50.615 ;
        RECT 56.535 46.655 57.175 1590.625 ;
        RECT 53.830 45.800 57.175 46.655 ;
        RECT 53.830 45.055 57.030 45.800 ;
        RECT 57.795 41.590 58.435 1591.885 ;
        RECT 55.165 40.595 58.435 41.590 ;
        RECT 55.165 39.990 58.365 40.595 ;
        RECT 59.095 36.640 59.735 1593.185 ;
        RECT 56.415 36.425 59.735 36.640 ;
        RECT 56.415 35.040 59.615 36.425 ;
        RECT 60.355 31.675 60.995 1594.445 ;
        RECT 57.725 30.075 60.995 31.675 ;
        RECT 60.355 29.870 60.995 30.075 ;
        RECT 61.655 26.690 62.295 1595.745 ;
        RECT 59.015 25.090 62.295 26.690 ;
        RECT 61.655 24.950 62.295 25.090 ;
        RECT 62.915 21.615 63.555 1597.005 ;
        RECT 60.220 20.715 63.555 21.615 ;
        RECT 60.220 20.015 63.420 20.715 ;
        RECT 64.215 16.650 64.855 1598.305 ;
        RECT 61.510 16.520 64.855 16.650 ;
        RECT 61.510 15.050 64.710 16.520 ;
        RECT 65.475 11.620 66.115 1599.565 ;
        RECT 62.780 10.020 66.115 11.620 ;
        RECT 65.475 9.945 66.115 10.020 ;
        RECT 66.775 6.720 67.415 1600.865 ;
        RECT 64.160 6.615 67.415 6.720 ;
        RECT 64.160 5.120 67.360 6.615 ;
        RECT 68.035 1.720 68.675 1602.125 ;
        RECT 69.335 6.720 69.975 1603.425 ;
        RECT 70.595 11.520 71.235 1604.685 ;
        RECT 70.595 9.920 73.985 11.520 ;
        RECT 70.595 9.670 71.235 9.920 ;
        RECT 69.335 6.620 72.605 6.720 ;
        RECT 69.405 5.120 72.605 6.620 ;
        RECT 97.660 6.570 99.530 6.610 ;
        RECT 96.245 4.970 99.530 6.570 ;
        RECT 97.660 1.935 99.530 4.970 ;
        RECT 68.035 0.120 71.355 1.720 ;
        RECT 68.035 0.000 68.675 0.120 ;
      LAYER met5 ;
        RECT 53.870 3868.380 57.310 3868.505 ;
        RECT 53.870 3866.780 214.605 3868.380 ;
        RECT 53.870 3866.665 57.310 3866.780 ;
        RECT 52.490 3863.380 55.930 3863.500 ;
        RECT 52.490 3861.780 217.910 3863.380 ;
        RECT 52.490 3861.660 55.930 3861.780 ;
        RECT 51.285 3858.380 54.725 3858.510 ;
        RECT 51.285 3856.780 214.605 3858.380 ;
        RECT 51.285 3856.670 54.725 3856.780 ;
        RECT 51.200 3763.380 54.640 3763.465 ;
        RECT 51.200 3761.780 214.605 3763.380 ;
        RECT 51.200 3761.625 54.640 3761.780 ;
        RECT 49.930 3758.380 53.370 3758.580 ;
        RECT 49.930 3756.780 217.910 3758.380 ;
        RECT 49.930 3756.740 53.370 3756.780 ;
        RECT 48.710 3753.380 52.150 3753.460 ;
        RECT 48.710 3751.780 214.605 3753.380 ;
        RECT 48.710 3751.620 52.150 3751.780 ;
        RECT 48.685 3658.380 52.125 3658.450 ;
        RECT 48.685 3656.780 214.605 3658.380 ;
        RECT 48.685 3656.610 52.125 3656.780 ;
        RECT 47.370 3653.380 50.810 3653.530 ;
        RECT 47.370 3651.780 217.910 3653.380 ;
        RECT 47.370 3651.690 50.810 3651.780 ;
        RECT 46.225 3648.380 49.665 3648.475 ;
        RECT 46.225 3646.780 214.605 3648.380 ;
        RECT 46.225 3646.635 49.665 3646.780 ;
        RECT 46.145 3553.380 49.585 3553.465 ;
        RECT 46.145 3551.780 214.605 3553.380 ;
        RECT 46.145 3551.625 49.585 3551.780 ;
        RECT 44.635 3548.380 48.075 3548.500 ;
        RECT 44.635 3546.780 217.905 3548.380 ;
        RECT 44.635 3546.660 48.075 3546.780 ;
        RECT 43.595 3543.380 47.035 3543.455 ;
        RECT 43.595 3541.780 214.605 3543.380 ;
        RECT 43.595 3541.615 47.035 3541.780 ;
        RECT 43.565 3102.270 47.005 3102.535 ;
        RECT 43.565 3100.695 214.605 3102.270 ;
        RECT 43.915 3100.670 214.605 3100.695 ;
        RECT 42.250 3097.270 45.690 3097.410 ;
        RECT 42.250 3095.670 217.905 3097.270 ;
        RECT 42.250 3095.570 45.690 3095.670 ;
        RECT 41.005 3092.270 44.445 3092.500 ;
        RECT 41.005 3090.670 214.605 3092.270 ;
        RECT 41.005 3090.660 44.445 3090.670 ;
        RECT 41.115 2937.270 44.555 2937.385 ;
        RECT 41.115 2935.670 214.605 2937.270 ;
        RECT 41.115 2935.545 44.555 2935.670 ;
        RECT 39.515 2932.270 42.955 2932.405 ;
        RECT 39.515 2930.670 217.905 2932.270 ;
        RECT 39.515 2930.565 42.955 2930.670 ;
        RECT 38.430 2927.270 41.870 2927.410 ;
        RECT 38.430 2925.670 214.605 2927.270 ;
        RECT 38.430 2925.570 41.870 2925.670 ;
        RECT 38.400 2772.270 41.840 2772.320 ;
        RECT 38.400 2770.670 214.605 2772.270 ;
        RECT 38.400 2770.480 41.840 2770.670 ;
        RECT 36.955 2767.270 40.395 2767.405 ;
        RECT 36.955 2765.670 217.905 2767.270 ;
        RECT 36.955 2765.565 40.395 2765.670 ;
        RECT 35.865 2762.270 39.305 2762.345 ;
        RECT 35.865 2760.670 214.605 2762.270 ;
        RECT 35.865 2760.505 39.305 2760.670 ;
        RECT 35.895 2607.270 39.335 2607.400 ;
        RECT 35.895 2605.670 214.605 2607.270 ;
        RECT 35.895 2605.560 39.335 2605.670 ;
        RECT 34.395 2602.270 37.835 2602.405 ;
        RECT 34.395 2600.670 217.905 2602.270 ;
        RECT 34.395 2600.565 37.835 2600.670 ;
        RECT 33.325 2597.270 36.765 2597.395 ;
        RECT 33.325 2595.670 214.605 2597.270 ;
        RECT 33.325 2595.555 36.765 2595.670 ;
        RECT 33.325 2288.345 36.765 2288.455 ;
        RECT 33.325 2286.745 214.605 2288.345 ;
        RECT 33.325 2286.615 36.765 2286.745 ;
        RECT 31.835 2283.345 35.275 2283.465 ;
        RECT 31.835 2281.745 217.905 2283.345 ;
        RECT 31.835 2281.625 35.275 2281.745 ;
        RECT 30.730 2278.345 34.170 2278.420 ;
        RECT 30.730 2276.745 214.605 2278.345 ;
        RECT 30.730 2276.580 34.170 2276.745 ;
        RECT 30.730 2119.270 34.170 2119.320 ;
        RECT 30.730 2117.670 214.605 2119.270 ;
        RECT 30.730 2117.480 34.170 2117.670 ;
        RECT 29.275 2114.270 32.715 2114.405 ;
        RECT 29.275 2112.670 217.905 2114.270 ;
        RECT 29.275 2112.565 32.715 2112.670 ;
        RECT 28.250 2109.270 31.690 2109.435 ;
        RECT 28.250 2107.670 214.605 2109.270 ;
        RECT 28.250 2107.595 31.690 2107.670 ;
        RECT 28.190 1954.270 31.630 1954.345 ;
        RECT 28.190 1952.670 214.605 1954.270 ;
        RECT 28.190 1952.505 31.630 1952.670 ;
        RECT 26.715 1949.270 30.155 1949.400 ;
        RECT 26.715 1947.670 217.905 1949.270 ;
        RECT 26.715 1947.560 30.155 1947.670 ;
        RECT 25.740 1944.270 29.180 1944.340 ;
        RECT 25.740 1942.670 214.605 1944.270 ;
        RECT 25.740 1942.500 29.180 1942.670 ;
        RECT 25.565 1787.840 29.005 1788.035 ;
        RECT 25.565 1786.240 214.605 1787.840 ;
        RECT 25.565 1786.195 29.005 1786.240 ;
        RECT 24.205 1782.840 27.645 1782.960 ;
        RECT 214.025 1782.840 217.905 1782.985 ;
        RECT 24.205 1781.385 217.905 1782.840 ;
        RECT 24.205 1781.240 217.745 1781.385 ;
        RECT 24.205 1781.120 27.645 1781.240 ;
        RECT 23.115 1777.840 26.555 1777.975 ;
        RECT 23.115 1776.240 214.605 1777.840 ;
        RECT 23.115 1776.135 26.555 1776.240 ;
        RECT 23.060 1622.985 26.500 1623.120 ;
        RECT 23.060 1621.385 214.605 1622.985 ;
        RECT 23.060 1621.280 26.500 1621.385 ;
        RECT 21.645 1617.985 25.085 1618.105 ;
        RECT 21.645 1616.385 217.905 1617.985 ;
        RECT 21.645 1616.265 25.085 1616.385 ;
        RECT 20.460 1612.985 23.900 1613.115 ;
        RECT 20.460 1611.385 214.605 1612.985 ;
        RECT 20.460 1611.275 23.900 1611.385 ;
        RECT 50.000 61.600 53.440 61.755 ;
        RECT 0.000 60.000 53.440 61.600 ;
        RECT 50.000 59.915 53.440 60.000 ;
        RECT 51.250 56.600 54.690 56.710 ;
        RECT 0.000 55.000 54.690 56.600 ;
        RECT 51.250 54.870 54.690 55.000 ;
        RECT 52.480 51.600 55.920 51.730 ;
        RECT 0.000 50.000 55.920 51.600 ;
        RECT 52.480 49.890 55.920 50.000 ;
        RECT 53.710 46.600 57.150 46.775 ;
        RECT 0.000 45.000 57.150 46.600 ;
        RECT 53.710 44.935 57.150 45.000 ;
        RECT 55.045 41.600 58.485 41.710 ;
        RECT 0.000 40.000 58.485 41.600 ;
        RECT 55.045 39.870 58.485 40.000 ;
        RECT 56.295 36.600 59.735 36.760 ;
        RECT 0.000 35.000 59.735 36.600 ;
        RECT 56.295 34.920 59.735 35.000 ;
        RECT 57.605 31.600 61.045 31.795 ;
        RECT 0.000 30.000 61.045 31.600 ;
        RECT 57.605 29.955 61.045 30.000 ;
        RECT 58.895 26.600 62.335 26.810 ;
        RECT 0.000 25.000 62.335 26.600 ;
        RECT 58.895 24.970 62.335 25.000 ;
        RECT 60.100 21.600 63.540 21.735 ;
        RECT 0.000 20.000 63.540 21.600 ;
        RECT 60.100 19.895 63.540 20.000 ;
        RECT 61.390 16.600 64.830 16.770 ;
        RECT 0.000 15.000 64.830 16.600 ;
        RECT 61.390 14.930 64.830 15.000 ;
        RECT 62.660 11.600 66.100 11.740 ;
        RECT 0.000 10.000 66.100 11.600 ;
        RECT 62.660 9.900 66.100 10.000 ;
        RECT 70.665 11.600 74.105 11.640 ;
        RECT 70.665 10.000 99.565 11.600 ;
        RECT 70.665 9.800 74.105 10.000 ;
        RECT 64.040 6.600 67.480 6.840 ;
        RECT 0.000 5.000 67.480 6.600 ;
        RECT 69.285 6.600 72.725 6.840 ;
        RECT 96.125 6.600 99.565 6.690 ;
        RECT 69.285 5.000 99.565 6.600 ;
        RECT 96.125 4.850 99.565 5.000 ;
        RECT 68.035 1.600 71.475 1.840 ;
        RECT 0.000 0.000 95.665 1.600 ;
  END
END analog_routes_right
END LIBRARY

