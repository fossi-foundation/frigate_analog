magic
tech sky130A
magscale 1 2
timestamp 1724444265
<< locali >>
rect 54 2797 12557 2922
<< metal1 >>
rect -186 2414 -180 2466
rect -128 2465 -122 2466
rect -128 2415 22 2465
rect 4232 2420 4238 2472
rect 4290 2471 4296 2472
rect 4290 2421 4550 2471
rect 4290 2420 4296 2421
rect 8766 2420 8772 2472
rect 8824 2471 8830 2472
rect 8824 2421 9062 2471
rect 8824 2420 8830 2421
rect -128 2414 -122 2415
rect -11 2037 335 2044
rect -11 1891 -2 2037
rect 324 1891 335 2037
rect 4505 2037 4851 2044
rect 4505 1891 4514 2037
rect 4840 1948 4851 2037
rect 9021 2037 9367 2044
rect 4840 1891 4857 1948
rect 9021 1891 9030 2037
rect 9356 1948 9367 2037
rect 9356 1891 9373 1948
rect -11 886 12565 1038
<< via1 >>
rect -180 2414 -128 2466
rect 2639 2461 3442 2548
rect 4238 2420 4290 2472
rect 7155 2461 7958 2548
rect 8772 2420 8824 2472
rect 11671 2461 12474 2548
rect -2 1891 324 2037
rect 4514 1891 4840 2037
rect 9030 1891 9356 2037
<< metal2 >>
rect 2622 2591 3465 2605
rect 2622 2565 2639 2591
rect -180 2466 -128 2472
rect 2625 2461 2639 2565
rect 3439 2569 3465 2591
rect 7138 2591 7981 2605
rect 3439 2548 3468 2569
rect 7138 2565 7155 2591
rect 3442 2461 3468 2548
rect 2625 2446 3468 2461
rect 4238 2472 4290 2478
rect 7141 2461 7155 2565
rect 7955 2569 7981 2591
rect 11654 2591 12497 2605
rect 7955 2548 7984 2569
rect 11654 2565 11671 2591
rect 7958 2461 7984 2548
rect 7141 2446 7984 2461
rect 8772 2472 8824 2478
rect 4238 2414 4290 2420
rect 11657 2461 11671 2565
rect 12471 2569 12497 2591
rect 12471 2548 12500 2569
rect 12474 2461 12500 2548
rect 11657 2446 12500 2461
rect 8772 2414 8824 2420
rect -180 2408 -128 2414
rect -179 896 -129 2408
rect -11 2037 335 2044
rect -11 1884 -2 2037
rect 324 1884 335 2037
rect -11 1879 335 1884
rect 4239 892 4289 2414
rect 4505 2037 4851 2044
rect 4505 1884 4514 2037
rect 4840 1884 4851 2037
rect 4505 1879 4851 1884
rect 8773 884 8823 2414
rect 9021 2037 9367 2044
rect 9021 1884 9030 2037
rect 9356 1884 9367 2037
rect 9021 1879 9367 1884
<< via2 >>
rect 942 4714 1887 4854
rect 5458 4714 6403 4854
rect 9974 4714 10919 4854
rect 742 3245 1687 3385
rect 5258 3245 6203 3385
rect 9774 3245 10719 3385
rect 2639 2548 3439 2591
rect 2639 2461 3439 2548
rect 7155 2548 7955 2591
rect 7155 2461 7955 2548
rect 11671 2548 12471 2591
rect 11671 2461 12471 2548
rect -2 1891 324 2037
rect -2 1884 324 1891
rect 4514 1891 4840 2037
rect 4514 1884 4840 1891
rect 9030 1891 9356 2037
rect 9030 1884 9356 1891
<< metal3 >>
rect -10 4854 12538 4884
rect -10 4714 942 4854
rect 1887 4714 5458 4854
rect 6403 4714 9974 4854
rect 10919 4714 12538 4854
rect -10 4705 12538 4714
rect -13 3385 12535 3407
rect -13 3245 742 3385
rect 1687 3245 5258 3385
rect 6203 3245 9774 3385
rect 10719 3245 12535 3385
rect -13 3228 12535 3245
rect 20 2591 12599 2606
rect 20 2461 2639 2591
rect 3439 2461 7155 2591
rect 7955 2461 11671 2591
rect 12471 2461 12599 2591
rect 20 2442 12599 2461
rect -17 2037 12580 2049
rect -17 1884 -2 2037
rect 324 1884 4514 2037
rect 4840 1884 9030 2037
rect 9356 1884 12580 2037
rect -17 1875 12580 1884
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_1 ../ip/sky130_ef_ip__analog_switches/mag
array 0 2 4516 0 0 -4247
timestamp 1724439637
transform 1 0 0 0 -1 4529
box -4 -600 3538 3648
<< end >>
