magic
tech sky130A
magscale 1 2
timestamp 1563080108
<< checkpaint >>
rect -1260 -1260 39379 503137
<< metal3 >>
rect 242 490293 942 490325
rect 242 490229 281 490293
rect 345 490229 361 490293
rect 425 490229 441 490293
rect 505 490229 521 490293
rect 585 490229 601 490293
rect 665 490229 681 490293
rect 745 490229 761 490293
rect 825 490229 841 490293
rect 905 490229 942 490293
rect 242 490197 942 490229
rect 242 469293 942 469325
rect 242 469229 281 469293
rect 345 469229 361 469293
rect 425 469229 441 469293
rect 505 469229 521 469293
rect 585 469229 601 469293
rect 665 469229 681 469293
rect 745 469229 761 469293
rect 825 469229 841 469293
rect 905 469229 942 469293
rect 242 469197 942 469229
rect 242 448293 942 448325
rect 242 448229 281 448293
rect 345 448229 361 448293
rect 425 448229 441 448293
rect 505 448229 521 448293
rect 585 448229 601 448293
rect 665 448229 681 448293
rect 745 448229 761 448293
rect 825 448229 841 448293
rect 905 448229 942 448293
rect 242 448197 942 448229
rect 242 427293 942 427325
rect 242 427229 281 427293
rect 345 427229 361 427293
rect 425 427229 441 427293
rect 505 427229 521 427293
rect 585 427229 601 427293
rect 665 427229 681 427293
rect 745 427229 761 427293
rect 825 427229 841 427293
rect 905 427229 942 427293
rect 242 427197 942 427229
rect 242 296547 942 296555
rect 0 296523 942 296547
rect 0 296459 281 296523
rect 345 296459 361 296523
rect 425 296459 441 296523
rect 505 296459 521 296523
rect 585 296459 601 296523
rect 665 296459 681 296523
rect 745 296459 761 296523
rect 825 296459 841 296523
rect 905 296459 942 296523
rect 0 296427 942 296459
rect 242 263547 942 263555
rect 0 263523 942 263547
rect 0 263459 281 263523
rect 345 263459 361 263523
rect 425 263459 441 263523
rect 505 263459 521 263523
rect 585 263459 601 263523
rect 665 263459 681 263523
rect 745 263459 761 263523
rect 825 263459 841 263523
rect 905 263459 942 263523
rect 0 263427 942 263459
rect 242 230547 942 230555
rect 0 230523 942 230547
rect 0 230459 281 230523
rect 345 230459 361 230523
rect 425 230459 441 230523
rect 505 230459 521 230523
rect 585 230459 601 230523
rect 665 230459 681 230523
rect 745 230459 761 230523
rect 825 230459 841 230523
rect 905 230459 942 230523
rect 0 230427 942 230459
rect 242 197547 942 197555
rect 0 197523 942 197547
rect 0 197459 281 197523
rect 345 197459 361 197523
rect 425 197459 441 197523
rect 505 197459 521 197523
rect 585 197459 601 197523
rect 665 197459 681 197523
rect 745 197459 761 197523
rect 825 197459 841 197523
rect 905 197459 942 197523
rect 0 197427 942 197459
rect 571 170411 871 170431
rect 571 170402 609 170411
rect 263 170002 609 170402
rect 571 169627 609 170002
rect 833 169627 871 170411
rect 571 169605 871 169627
rect 242 160100 942 160132
rect 242 160036 281 160100
rect 345 160036 361 160100
rect 425 160036 441 160100
rect 505 160036 521 160100
rect 585 160036 601 160100
rect 665 160036 681 160100
rect 745 160036 761 160100
rect 825 160036 841 160100
rect 905 160036 942 160100
rect 242 160004 942 160036
rect 242 99947 942 99955
rect 241 99923 942 99947
rect 241 99859 281 99923
rect 345 99859 361 99923
rect 425 99859 441 99923
rect 505 99859 521 99923
rect 585 99859 601 99923
rect 665 99859 681 99923
rect 745 99859 761 99923
rect 825 99859 841 99923
rect 905 99859 942 99923
rect 241 99827 942 99859
rect 242 66947 942 66955
rect 0 66923 942 66947
rect 0 66859 281 66923
rect 345 66859 361 66923
rect 425 66859 441 66923
rect 505 66859 521 66923
rect 585 66859 601 66923
rect 665 66859 681 66923
rect 745 66859 761 66923
rect 825 66859 841 66923
rect 905 66859 942 66923
rect 0 66827 942 66859
rect 242 34204 942 34212
rect 0 34180 942 34204
rect 0 34116 281 34180
rect 345 34116 361 34180
rect 425 34116 441 34180
rect 505 34116 521 34180
rect 585 34116 601 34180
rect 665 34116 681 34180
rect 745 34116 761 34180
rect 825 34116 841 34180
rect 905 34116 942 34180
rect 0 34084 942 34116
rect 242 1204 942 1212
rect 0 1180 942 1204
rect 0 1116 281 1180
rect 345 1116 361 1180
rect 425 1116 441 1180
rect 505 1116 521 1180
rect 585 1116 601 1180
rect 665 1116 681 1180
rect 745 1116 761 1180
rect 825 1116 841 1180
rect 905 1116 942 1180
rect 0 1084 942 1116
<< via3 >>
rect 281 490229 345 490293
rect 361 490229 425 490293
rect 441 490229 505 490293
rect 521 490229 585 490293
rect 601 490229 665 490293
rect 681 490229 745 490293
rect 761 490229 825 490293
rect 841 490229 905 490293
rect 281 469229 345 469293
rect 361 469229 425 469293
rect 441 469229 505 469293
rect 521 469229 585 469293
rect 601 469229 665 469293
rect 681 469229 745 469293
rect 761 469229 825 469293
rect 841 469229 905 469293
rect 281 448229 345 448293
rect 361 448229 425 448293
rect 441 448229 505 448293
rect 521 448229 585 448293
rect 601 448229 665 448293
rect 681 448229 745 448293
rect 761 448229 825 448293
rect 841 448229 905 448293
rect 281 427229 345 427293
rect 361 427229 425 427293
rect 441 427229 505 427293
rect 521 427229 585 427293
rect 601 427229 665 427293
rect 681 427229 745 427293
rect 761 427229 825 427293
rect 841 427229 905 427293
rect 281 296459 345 296523
rect 361 296459 425 296523
rect 441 296459 505 296523
rect 521 296459 585 296523
rect 601 296459 665 296523
rect 681 296459 745 296523
rect 761 296459 825 296523
rect 841 296459 905 296523
rect 281 263459 345 263523
rect 361 263459 425 263523
rect 441 263459 505 263523
rect 521 263459 585 263523
rect 601 263459 665 263523
rect 681 263459 745 263523
rect 761 263459 825 263523
rect 841 263459 905 263523
rect 281 230459 345 230523
rect 361 230459 425 230523
rect 441 230459 505 230523
rect 521 230459 585 230523
rect 601 230459 665 230523
rect 681 230459 745 230523
rect 761 230459 825 230523
rect 841 230459 905 230523
rect 281 197459 345 197523
rect 361 197459 425 197523
rect 441 197459 505 197523
rect 521 197459 585 197523
rect 601 197459 665 197523
rect 681 197459 745 197523
rect 761 197459 825 197523
rect 841 197459 905 197523
rect 609 169627 833 170411
rect 281 160036 345 160100
rect 361 160036 425 160100
rect 441 160036 505 160100
rect 521 160036 585 160100
rect 601 160036 665 160100
rect 681 160036 745 160100
rect 761 160036 825 160100
rect 841 160036 905 160100
rect 281 99859 345 99923
rect 361 99859 425 99923
rect 441 99859 505 99923
rect 521 99859 585 99923
rect 601 99859 665 99923
rect 681 99859 745 99923
rect 761 99859 825 99923
rect 841 99859 905 99923
rect 281 66859 345 66923
rect 361 66859 425 66923
rect 441 66859 505 66923
rect 521 66859 585 66923
rect 601 66859 665 66923
rect 681 66859 745 66923
rect 761 66859 825 66923
rect 841 66859 905 66923
rect 281 34116 345 34180
rect 361 34116 425 34180
rect 441 34116 505 34180
rect 521 34116 585 34180
rect 601 34116 665 34180
rect 681 34116 745 34180
rect 761 34116 825 34180
rect 841 34116 905 34180
rect 281 1116 345 1180
rect 361 1116 425 1180
rect 441 1116 505 1180
rect 521 1116 585 1180
rect 601 1116 665 1180
rect 681 1116 745 1180
rect 761 1116 825 1180
rect 841 1116 905 1180
<< metal4 >>
rect 31327 491433 31455 501877
rect 30814 491391 31455 491433
rect 30814 491155 30856 491391
rect 31092 491155 31176 491391
rect 31412 491155 31455 491391
rect 30814 491113 31455 491155
rect 31327 491112 31455 491113
rect 31587 490433 31715 501877
rect 452 490391 948 490433
rect 452 490325 586 490391
rect 242 490293 586 490325
rect 822 490293 948 490391
rect 242 490229 281 490293
rect 345 490229 361 490293
rect 425 490229 441 490293
rect 505 490229 521 490293
rect 585 490229 586 490293
rect 825 490229 841 490293
rect 905 490229 948 490293
rect 242 490197 586 490229
rect 452 490155 586 490197
rect 822 490155 948 490229
rect 452 490113 948 490155
rect 31075 490391 31715 490433
rect 31075 490155 31117 490391
rect 31353 490155 31437 490391
rect 31673 490155 31715 490391
rect 31075 490113 31715 490155
rect 31839 489433 31967 501877
rect 31327 489391 31967 489433
rect 31327 489155 31369 489391
rect 31605 489155 31689 489391
rect 31925 489155 31967 489391
rect 31327 489113 31967 489155
rect 31839 470433 31967 489113
rect 31326 470391 31967 470433
rect 31326 470155 31368 470391
rect 31604 470155 31688 470391
rect 31924 470155 31967 470391
rect 31326 470113 31967 470155
rect 31839 470111 31967 470113
rect 32099 469433 32227 501877
rect 452 469391 948 469433
rect 452 469325 586 469391
rect 242 469293 586 469325
rect 822 469293 948 469391
rect 242 469229 281 469293
rect 345 469229 361 469293
rect 425 469229 441 469293
rect 505 469229 521 469293
rect 585 469229 586 469293
rect 825 469229 841 469293
rect 905 469229 948 469293
rect 242 469197 586 469229
rect 452 469155 586 469197
rect 822 469155 948 469229
rect 452 469113 948 469155
rect 31588 469391 32228 469433
rect 31588 469155 31630 469391
rect 31866 469155 31950 469391
rect 32186 469155 32228 469391
rect 31588 469113 32228 469155
rect 32351 468433 32479 501877
rect 31839 468391 32479 468433
rect 31839 468155 31881 468391
rect 32117 468155 32201 468391
rect 32437 468155 32479 468391
rect 31839 468113 32479 468155
rect 32351 449434 32479 468113
rect 31839 449392 32479 449434
rect 31839 449156 31881 449392
rect 32117 449156 32201 449392
rect 32437 449156 32479 449392
rect 31839 449114 32479 449156
rect 32351 449112 32479 449114
rect 32611 448433 32739 501877
rect 452 448391 948 448433
rect 452 448325 586 448391
rect 242 448293 586 448325
rect 822 448293 948 448391
rect 242 448229 281 448293
rect 345 448229 361 448293
rect 425 448229 441 448293
rect 505 448229 521 448293
rect 585 448229 586 448293
rect 825 448229 841 448293
rect 905 448229 948 448293
rect 242 448197 586 448229
rect 452 448155 586 448197
rect 822 448155 948 448229
rect 452 448113 948 448155
rect 32099 448391 32739 448433
rect 32099 448155 32141 448391
rect 32377 448155 32461 448391
rect 32697 448155 32739 448391
rect 32099 448113 32739 448155
rect 32863 447432 32991 501877
rect 32350 447390 32991 447432
rect 32350 447154 32392 447390
rect 32628 447154 32712 447390
rect 32948 447154 32991 447390
rect 32350 447112 32991 447154
rect 32863 428433 32991 447112
rect 32351 428391 32991 428433
rect 32351 428155 32393 428391
rect 32629 428155 32713 428391
rect 32949 428155 32991 428391
rect 32351 428113 32991 428155
rect 32863 428103 32991 428113
rect 33123 427433 33251 501877
rect 452 427391 948 427433
rect 452 427325 586 427391
rect 242 427293 586 427325
rect 822 427293 948 427391
rect 242 427229 281 427293
rect 345 427229 361 427293
rect 425 427229 441 427293
rect 505 427229 521 427293
rect 585 427229 586 427293
rect 825 427229 841 427293
rect 905 427229 948 427293
rect 242 427197 586 427229
rect 452 427155 586 427197
rect 822 427155 948 427229
rect 452 427113 948 427155
rect 32612 427391 33252 427433
rect 32612 427155 32654 427391
rect 32890 427155 32974 427391
rect 33210 427155 33252 427391
rect 32612 427113 33252 427155
rect 33375 426435 33503 501877
rect 32864 426393 33504 426435
rect 32864 426157 32906 426393
rect 33142 426157 33226 426393
rect 33462 426157 33504 426393
rect 32864 426115 33504 426157
rect 33375 297661 33503 426115
rect 32863 297619 33503 297661
rect 32863 297383 32905 297619
rect 33141 297383 33225 297619
rect 33461 297383 33503 297619
rect 32863 297341 33503 297383
rect 33635 296665 33763 501877
rect 452 296621 948 296664
rect 452 296555 586 296621
rect 242 296523 586 296555
rect 822 296523 948 296621
rect 242 296459 281 296523
rect 345 296459 361 296523
rect 425 296459 441 296523
rect 505 296459 521 296523
rect 585 296459 586 296523
rect 825 296459 841 296523
rect 905 296459 948 296523
rect 242 296427 586 296459
rect 452 296385 586 296427
rect 822 296385 948 296459
rect 452 296343 948 296385
rect 33123 296623 33763 296665
rect 33123 296387 33165 296623
rect 33401 296387 33485 296623
rect 33721 296387 33763 296623
rect 33123 296345 33763 296387
rect 33887 295661 34015 501877
rect 33376 295619 34016 295661
rect 33376 295383 33418 295619
rect 33654 295383 33738 295619
rect 33974 295383 34016 295619
rect 33376 295341 34016 295383
rect 33887 264660 34015 295341
rect 33376 264618 34016 264660
rect 33376 264382 33418 264618
rect 33654 264382 33738 264618
rect 33974 264382 34016 264618
rect 33376 264340 34016 264382
rect 33887 264336 34015 264340
rect 452 263621 948 263663
rect 34147 263659 34275 501877
rect 452 263555 586 263621
rect 242 263523 586 263555
rect 822 263523 948 263621
rect 242 263459 281 263523
rect 345 263459 361 263523
rect 425 263459 441 263523
rect 505 263459 521 263523
rect 585 263459 586 263523
rect 825 263459 841 263523
rect 905 263459 948 263523
rect 242 263427 586 263459
rect 452 263385 586 263427
rect 822 263385 948 263459
rect 452 263343 948 263385
rect 33635 263617 34275 263659
rect 33635 263381 33677 263617
rect 33913 263381 33997 263617
rect 34233 263381 34275 263617
rect 33635 263339 34275 263381
rect 34399 262661 34527 501877
rect 33887 262619 34527 262661
rect 33887 262383 33929 262619
rect 34165 262383 34249 262619
rect 34485 262383 34527 262619
rect 33887 262341 34527 262383
rect 34399 231685 34527 262341
rect 33888 231643 34528 231685
rect 33888 231407 33930 231643
rect 34166 231407 34250 231643
rect 34486 231407 34528 231643
rect 33888 231365 34528 231407
rect 34399 231361 34527 231365
rect 34659 230687 34787 501877
rect 452 230621 948 230663
rect 452 230555 586 230621
rect 242 230523 586 230555
rect 822 230523 948 230621
rect 242 230459 281 230523
rect 345 230459 361 230523
rect 425 230459 441 230523
rect 505 230459 521 230523
rect 585 230459 586 230523
rect 825 230459 841 230523
rect 905 230459 948 230523
rect 242 230427 586 230459
rect 452 230385 586 230427
rect 822 230385 948 230459
rect 452 230343 948 230385
rect 34147 230645 34787 230687
rect 34147 230409 34189 230645
rect 34425 230409 34509 230645
rect 34745 230409 34787 230645
rect 34147 230367 34787 230409
rect 34911 229688 35039 501877
rect 34400 229646 35040 229688
rect 34400 229410 34442 229646
rect 34678 229410 34762 229646
rect 34998 229410 35040 229646
rect 34400 229368 35040 229410
rect 34911 198660 35039 229368
rect 34399 198618 35039 198660
rect 34399 198382 34441 198618
rect 34677 198382 34761 198618
rect 34997 198382 35039 198618
rect 34399 198340 35039 198382
rect 452 197621 948 197663
rect 35171 197662 35299 501877
rect 452 197555 586 197621
rect 242 197523 586 197555
rect 822 197523 948 197621
rect 242 197459 281 197523
rect 345 197459 361 197523
rect 425 197459 441 197523
rect 505 197459 521 197523
rect 585 197459 586 197523
rect 825 197459 841 197523
rect 905 197459 948 197523
rect 242 197427 586 197459
rect 452 197385 586 197427
rect 822 197385 948 197459
rect 452 197343 948 197385
rect 34659 197620 35299 197662
rect 34659 197384 34701 197620
rect 34937 197384 35021 197620
rect 35257 197384 35299 197620
rect 34659 197342 35299 197384
rect 35423 196661 35551 501877
rect 34913 196619 35553 196661
rect 34913 196383 34955 196619
rect 35191 196383 35275 196619
rect 35511 196383 35553 196619
rect 34913 196341 35553 196383
rect 571 170411 871 170431
rect 571 169627 609 170411
rect 833 169627 871 170411
rect 571 169605 871 169627
rect 645 160240 797 169605
rect 35423 161241 35551 196341
rect 34911 161199 35551 161241
rect 34911 160963 34953 161199
rect 35189 160963 35273 161199
rect 35509 160963 35551 161199
rect 34911 160921 35551 160963
rect 35423 160919 35551 160921
rect 35683 160240 35811 501877
rect 452 160198 948 160240
rect 452 160132 586 160198
rect 242 160100 586 160132
rect 822 160100 948 160198
rect 242 160036 281 160100
rect 345 160036 361 160100
rect 425 160036 441 160100
rect 505 160036 521 160100
rect 585 160036 586 160100
rect 825 160036 841 160100
rect 905 160036 948 160100
rect 242 160004 586 160036
rect 452 159962 586 160004
rect 822 159962 948 160036
rect 452 159920 948 159962
rect 35171 160198 35811 160240
rect 35171 159962 35213 160198
rect 35449 159962 35533 160198
rect 35769 159962 35811 160198
rect 35171 159920 35811 159962
rect 35935 159241 36063 501877
rect 35422 159199 36063 159241
rect 35422 158963 35464 159199
rect 35700 158963 35784 159199
rect 36020 158963 36063 159199
rect 35422 158921 36063 158963
rect 35935 101060 36063 158921
rect 35423 101018 36063 101060
rect 35423 100782 35465 101018
rect 35701 100782 35785 101018
rect 36021 100782 36063 101018
rect 35423 100740 36063 100782
rect 452 100021 948 100063
rect 36195 100062 36323 501877
rect 452 99955 586 100021
rect 242 99923 586 99955
rect 822 99923 948 100021
rect 242 99859 281 99923
rect 345 99859 361 99923
rect 425 99859 441 99923
rect 505 99859 521 99923
rect 585 99859 586 99923
rect 825 99859 841 99923
rect 905 99859 948 99923
rect 242 99827 586 99859
rect 452 99785 586 99827
rect 822 99785 948 99859
rect 452 99743 948 99785
rect 35685 100020 36325 100062
rect 35685 99784 35727 100020
rect 35963 99784 36047 100020
rect 36283 99784 36325 100020
rect 35685 99742 36325 99784
rect 36447 99062 36575 501877
rect 35935 99020 36575 99062
rect 35935 98784 35977 99020
rect 36213 98784 36297 99020
rect 36533 98784 36575 99020
rect 35935 98742 36575 98784
rect 36447 68059 36575 98742
rect 35933 68017 36575 68059
rect 35933 67781 35975 68017
rect 36211 67781 36295 68017
rect 36531 67781 36575 68017
rect 35933 67741 36575 67781
rect 35933 67739 36573 67741
rect 452 67021 948 67063
rect 36707 67059 36835 501877
rect 452 66955 586 67021
rect 242 66923 586 66955
rect 822 66923 948 67021
rect 242 66859 281 66923
rect 345 66859 361 66923
rect 425 66859 441 66923
rect 505 66859 521 66923
rect 585 66859 586 66923
rect 825 66859 841 66923
rect 905 66859 948 66923
rect 242 66827 586 66859
rect 452 66785 586 66827
rect 822 66785 948 66859
rect 452 66743 948 66785
rect 36195 67017 36835 67059
rect 36195 66781 36237 67017
rect 36473 66781 36557 67017
rect 36793 66781 36835 67017
rect 36195 66739 36835 66781
rect 36959 66059 37087 501877
rect 36447 66017 37087 66059
rect 36447 65781 36489 66017
rect 36725 65781 36809 66017
rect 37045 65781 37087 66017
rect 36447 65739 37087 65781
rect 36959 35321 37087 65739
rect 36447 35279 37087 35321
rect 36447 35043 36489 35279
rect 36725 35043 36809 35279
rect 37045 35043 37087 35279
rect 36447 35001 37087 35043
rect 452 34278 948 34320
rect 37219 34315 37347 501877
rect 452 34212 586 34278
rect 242 34180 586 34212
rect 822 34180 948 34278
rect 242 34116 281 34180
rect 345 34116 361 34180
rect 425 34116 441 34180
rect 505 34116 521 34180
rect 585 34116 586 34180
rect 825 34116 841 34180
rect 905 34116 948 34180
rect 242 34084 586 34116
rect 452 34042 586 34084
rect 822 34042 948 34116
rect 452 34000 948 34042
rect 36707 34273 37347 34315
rect 36707 34037 36749 34273
rect 36985 34037 37069 34273
rect 37305 34037 37347 34273
rect 36707 33995 37347 34037
rect 37471 33321 37599 501877
rect 36960 33279 37600 33321
rect 36960 33043 37002 33279
rect 37238 33043 37322 33279
rect 37558 33043 37600 33279
rect 36960 33001 37600 33043
rect 37471 2315 37599 33001
rect 36935 2273 37599 2315
rect 36935 2037 36977 2273
rect 37213 2037 37297 2273
rect 37533 2037 37599 2273
rect 36935 1995 37599 2037
rect 37471 1987 37599 1995
rect 452 1278 948 1320
rect 37731 1319 37859 501877
rect 452 1212 586 1278
rect 242 1180 586 1212
rect 822 1180 948 1278
rect 242 1116 281 1180
rect 345 1116 361 1180
rect 425 1116 441 1180
rect 505 1116 521 1180
rect 585 1116 586 1180
rect 825 1116 841 1180
rect 905 1116 948 1180
rect 242 1084 586 1116
rect 452 1042 586 1084
rect 822 1042 948 1116
rect 452 1000 948 1042
rect 37219 1277 37859 1319
rect 37219 1041 37261 1277
rect 37497 1041 37581 1277
rect 37817 1041 37859 1277
rect 37219 999 37859 1041
rect 37991 344 38119 501877
rect 37455 302 38119 344
rect 37455 66 37497 302
rect 37733 66 37817 302
rect 38053 66 38119 302
rect 37455 24 38119 66
rect 37991 0 38119 24
<< via4 >>
rect 30856 491155 31092 491391
rect 31176 491155 31412 491391
rect 586 490293 822 490391
rect 586 490229 601 490293
rect 601 490229 665 490293
rect 665 490229 681 490293
rect 681 490229 745 490293
rect 745 490229 761 490293
rect 761 490229 822 490293
rect 586 490155 822 490229
rect 31117 490155 31353 490391
rect 31437 490155 31673 490391
rect 31369 489155 31605 489391
rect 31689 489155 31925 489391
rect 31368 470155 31604 470391
rect 31688 470155 31924 470391
rect 586 469293 822 469391
rect 586 469229 601 469293
rect 601 469229 665 469293
rect 665 469229 681 469293
rect 681 469229 745 469293
rect 745 469229 761 469293
rect 761 469229 822 469293
rect 586 469155 822 469229
rect 31630 469155 31866 469391
rect 31950 469155 32186 469391
rect 31881 468155 32117 468391
rect 32201 468155 32437 468391
rect 31881 449156 32117 449392
rect 32201 449156 32437 449392
rect 586 448293 822 448391
rect 586 448229 601 448293
rect 601 448229 665 448293
rect 665 448229 681 448293
rect 681 448229 745 448293
rect 745 448229 761 448293
rect 761 448229 822 448293
rect 586 448155 822 448229
rect 32141 448155 32377 448391
rect 32461 448155 32697 448391
rect 32392 447154 32628 447390
rect 32712 447154 32948 447390
rect 32393 428155 32629 428391
rect 32713 428155 32949 428391
rect 586 427293 822 427391
rect 586 427229 601 427293
rect 601 427229 665 427293
rect 665 427229 681 427293
rect 681 427229 745 427293
rect 745 427229 761 427293
rect 761 427229 822 427293
rect 586 427155 822 427229
rect 32654 427155 32890 427391
rect 32974 427155 33210 427391
rect 32906 426157 33142 426393
rect 33226 426157 33462 426393
rect 32905 297383 33141 297619
rect 33225 297383 33461 297619
rect 586 296523 822 296621
rect 586 296459 601 296523
rect 601 296459 665 296523
rect 665 296459 681 296523
rect 681 296459 745 296523
rect 745 296459 761 296523
rect 761 296459 822 296523
rect 586 296385 822 296459
rect 33165 296387 33401 296623
rect 33485 296387 33721 296623
rect 33418 295383 33654 295619
rect 33738 295383 33974 295619
rect 33418 264382 33654 264618
rect 33738 264382 33974 264618
rect 586 263523 822 263621
rect 586 263459 601 263523
rect 601 263459 665 263523
rect 665 263459 681 263523
rect 681 263459 745 263523
rect 745 263459 761 263523
rect 761 263459 822 263523
rect 586 263385 822 263459
rect 33677 263381 33913 263617
rect 33997 263381 34233 263617
rect 33929 262383 34165 262619
rect 34249 262383 34485 262619
rect 33930 231407 34166 231643
rect 34250 231407 34486 231643
rect 586 230523 822 230621
rect 586 230459 601 230523
rect 601 230459 665 230523
rect 665 230459 681 230523
rect 681 230459 745 230523
rect 745 230459 761 230523
rect 761 230459 822 230523
rect 586 230385 822 230459
rect 34189 230409 34425 230645
rect 34509 230409 34745 230645
rect 34442 229410 34678 229646
rect 34762 229410 34998 229646
rect 34441 198382 34677 198618
rect 34761 198382 34997 198618
rect 586 197523 822 197621
rect 586 197459 601 197523
rect 601 197459 665 197523
rect 665 197459 681 197523
rect 681 197459 745 197523
rect 745 197459 761 197523
rect 761 197459 822 197523
rect 586 197385 822 197459
rect 34701 197384 34937 197620
rect 35021 197384 35257 197620
rect 34955 196383 35191 196619
rect 35275 196383 35511 196619
rect 34953 160963 35189 161199
rect 35273 160963 35509 161199
rect 586 160100 822 160198
rect 586 160036 601 160100
rect 601 160036 665 160100
rect 665 160036 681 160100
rect 681 160036 745 160100
rect 745 160036 761 160100
rect 761 160036 822 160100
rect 586 159962 822 160036
rect 35213 159962 35449 160198
rect 35533 159962 35769 160198
rect 35464 158963 35700 159199
rect 35784 158963 36020 159199
rect 35465 100782 35701 101018
rect 35785 100782 36021 101018
rect 586 99923 822 100021
rect 586 99859 601 99923
rect 601 99859 665 99923
rect 665 99859 681 99923
rect 681 99859 745 99923
rect 745 99859 761 99923
rect 761 99859 822 99923
rect 586 99785 822 99859
rect 35727 99784 35963 100020
rect 36047 99784 36283 100020
rect 35977 98784 36213 99020
rect 36297 98784 36533 99020
rect 35975 67781 36211 68017
rect 36295 67781 36531 68017
rect 586 66923 822 67021
rect 586 66859 601 66923
rect 601 66859 665 66923
rect 665 66859 681 66923
rect 681 66859 745 66923
rect 745 66859 761 66923
rect 761 66859 822 66923
rect 586 66785 822 66859
rect 36237 66781 36473 67017
rect 36557 66781 36793 67017
rect 36489 65781 36725 66017
rect 36809 65781 37045 66017
rect 36489 35043 36725 35279
rect 36809 35043 37045 35279
rect 586 34180 822 34278
rect 586 34116 601 34180
rect 601 34116 665 34180
rect 665 34116 681 34180
rect 681 34116 745 34180
rect 745 34116 761 34180
rect 761 34116 822 34180
rect 586 34042 822 34116
rect 36749 34037 36985 34273
rect 37069 34037 37305 34273
rect 37002 33043 37238 33279
rect 37322 33043 37558 33279
rect 36977 2037 37213 2273
rect 37297 2037 37533 2273
rect 586 1180 822 1278
rect 586 1116 601 1180
rect 601 1116 665 1180
rect 665 1116 681 1180
rect 681 1116 745 1180
rect 745 1116 761 1180
rect 761 1116 822 1180
rect 586 1042 822 1116
rect 37261 1041 37497 1277
rect 37581 1041 37817 1277
rect 37497 66 37733 302
rect 37817 66 38053 302
<< metal5 >>
rect 30790 491433 31478 491457
rect 924 491391 31491 491433
rect 924 491155 30856 491391
rect 31092 491155 31176 491391
rect 31412 491155 31491 491391
rect 924 491113 31491 491155
rect 30790 491089 31478 491113
rect 31051 490433 31739 490457
rect 452 490391 31739 490433
rect 452 490155 586 490391
rect 822 490155 31117 490391
rect 31353 490155 31437 490391
rect 31673 490155 31739 490391
rect 452 490113 31739 490155
rect 31051 490089 31739 490113
rect 31303 489433 31991 489457
rect 924 489391 31991 489433
rect 924 489155 31369 489391
rect 31605 489155 31689 489391
rect 31925 489155 31991 489391
rect 924 489113 31991 489155
rect 31303 489089 31991 489113
rect 31302 470433 31990 470457
rect 924 470391 32003 470433
rect 924 470155 31368 470391
rect 31604 470155 31688 470391
rect 31924 470155 32003 470391
rect 924 470113 32003 470155
rect 31302 470089 31990 470113
rect 31564 469433 32252 469457
rect 452 469391 32252 469433
rect 452 469155 586 469391
rect 822 469155 31630 469391
rect 31866 469155 31950 469391
rect 32186 469155 32252 469391
rect 452 469113 32252 469155
rect 31564 469089 32252 469113
rect 31815 468433 32503 468457
rect 924 468391 32503 468433
rect 924 468155 31881 468391
rect 32117 468155 32201 468391
rect 32437 468155 32503 468391
rect 924 468113 32503 468155
rect 31815 468089 32503 468113
rect 31815 449433 32503 449458
rect 924 449392 32515 449433
rect 924 449156 31881 449392
rect 32117 449156 32201 449392
rect 32437 449156 32515 449392
rect 924 449113 32515 449156
rect 31815 449090 32503 449113
rect 32075 448433 32763 448457
rect 452 448391 32763 448433
rect 452 448155 586 448391
rect 822 448155 32141 448391
rect 32377 448155 32461 448391
rect 32697 448155 32763 448391
rect 452 448113 32763 448155
rect 32075 448089 32763 448113
rect 32326 447433 33014 447456
rect 924 447390 33014 447433
rect 924 447154 32392 447390
rect 32628 447154 32712 447390
rect 32948 447154 33014 447390
rect 924 447113 33014 447154
rect 32326 447088 33014 447113
rect 32327 428433 33015 428457
rect 924 428391 33027 428433
rect 924 428155 32393 428391
rect 32629 428155 32713 428391
rect 32949 428155 33027 428391
rect 924 428113 33027 428155
rect 32327 428089 33015 428113
rect 32588 427433 33276 427457
rect 452 427391 33276 427433
rect 452 427155 586 427391
rect 822 427155 32654 427391
rect 32890 427155 32974 427391
rect 33210 427155 33276 427391
rect 452 427113 33276 427155
rect 32588 427089 33276 427113
rect 32840 426433 33528 426459
rect 924 426393 33528 426433
rect 924 426157 32906 426393
rect 33142 426157 33226 426393
rect 33462 426157 33528 426393
rect 924 426113 33528 426157
rect 32840 426091 33528 426113
rect 32839 297664 33527 297685
rect 924 297619 33539 297664
rect 924 297383 32905 297619
rect 33141 297383 33225 297619
rect 33461 297383 33539 297619
rect 924 297344 33539 297383
rect 32839 297317 33527 297344
rect 33099 296664 33787 296689
rect 452 296623 33787 296664
rect 452 296621 33165 296623
rect 452 296385 586 296621
rect 822 296387 33165 296621
rect 33401 296387 33485 296623
rect 33721 296387 33787 296623
rect 822 296385 33787 296387
rect 452 296344 33787 296385
rect 33099 296321 33787 296344
rect 33352 295664 34040 295685
rect 924 295619 34040 295664
rect 924 295383 33418 295619
rect 33654 295383 33738 295619
rect 33974 295383 34040 295619
rect 924 295344 34040 295383
rect 33352 295317 34040 295344
rect 33352 264663 34040 264684
rect 924 264618 34051 264663
rect 924 264382 33418 264618
rect 33654 264382 33738 264618
rect 33974 264382 34051 264618
rect 924 264343 34051 264382
rect 33352 264316 34040 264343
rect 33611 263663 34299 263683
rect 452 263621 34299 263663
rect 452 263385 586 263621
rect 822 263617 34299 263621
rect 822 263385 33677 263617
rect 452 263381 33677 263385
rect 33913 263381 33997 263617
rect 34233 263381 34299 263617
rect 452 263343 34299 263381
rect 33611 263315 34299 263343
rect 33863 262663 34551 262685
rect 924 262619 34551 262663
rect 924 262383 33929 262619
rect 34165 262383 34249 262619
rect 34485 262383 34551 262619
rect 924 262343 34551 262383
rect 33863 262317 34551 262343
rect 33864 231690 34552 231709
rect 924 231643 34563 231690
rect 924 231407 33930 231643
rect 34166 231407 34250 231643
rect 34486 231407 34563 231643
rect 924 231370 34563 231407
rect 33864 231341 34552 231370
rect 34123 230690 34811 230711
rect 603 230663 34811 230690
rect 452 230645 34811 230663
rect 452 230621 34189 230645
rect 452 230385 586 230621
rect 822 230409 34189 230621
rect 34425 230409 34509 230645
rect 34745 230409 34811 230645
rect 822 230385 34811 230409
rect 452 230370 34811 230385
rect 452 230343 1013 230370
rect 34123 230343 34811 230370
rect 34376 229690 35064 229712
rect 924 229646 35064 229690
rect 924 229410 34442 229646
rect 34678 229410 34762 229646
rect 34998 229410 35064 229646
rect 924 229370 35064 229410
rect 34376 229344 35064 229370
rect 34375 198663 35063 198684
rect 924 198618 35075 198663
rect 924 198382 34441 198618
rect 34677 198382 34761 198618
rect 34997 198382 35075 198618
rect 924 198343 35075 198382
rect 34375 198316 35063 198343
rect 34635 197663 35323 197686
rect 452 197621 35323 197663
rect 452 197385 586 197621
rect 822 197620 35323 197621
rect 822 197385 34701 197620
rect 452 197384 34701 197385
rect 34937 197384 35021 197620
rect 35257 197384 35323 197620
rect 452 197343 35323 197384
rect 34635 197318 35323 197343
rect 34889 196663 35577 196685
rect 924 196619 35577 196663
rect 924 196383 34955 196619
rect 35191 196383 35275 196619
rect 35511 196383 35577 196619
rect 924 196343 35577 196383
rect 34889 196317 35577 196343
rect 34887 161240 35575 161265
rect 924 161199 35587 161240
rect 924 160963 34953 161199
rect 35189 160963 35273 161199
rect 35509 160963 35587 161199
rect 924 160920 35587 160963
rect 34887 160897 35575 160920
rect 35147 160240 35835 160264
rect 452 160198 35835 160240
rect 452 159962 586 160198
rect 822 159962 35213 160198
rect 35449 159962 35533 160198
rect 35769 159962 35835 160198
rect 452 159920 35835 159962
rect 35147 159896 35835 159920
rect 35398 159240 36086 159265
rect 924 159199 36086 159240
rect 924 158963 35464 159199
rect 35700 158963 35784 159199
rect 36020 158963 36086 159199
rect 924 158920 36086 158963
rect 35398 158897 36086 158920
rect 35399 101063 36087 101084
rect 924 101018 36099 101063
rect 924 100782 35465 101018
rect 35701 100782 35785 101018
rect 36021 100782 36099 101018
rect 924 100743 36099 100782
rect 35399 100716 36087 100743
rect 35661 100063 36349 100086
rect 452 100021 36349 100063
rect 452 99785 586 100021
rect 822 100020 36349 100021
rect 822 99785 35727 100020
rect 452 99784 35727 99785
rect 35963 99784 36047 100020
rect 36283 99784 36349 100020
rect 452 99743 36349 99784
rect 35661 99718 36349 99743
rect 35911 99063 36599 99086
rect 924 99020 36599 99063
rect 924 98784 35977 99020
rect 36213 98784 36297 99020
rect 36533 98784 36599 99020
rect 924 98743 36599 98784
rect 35911 98718 36599 98743
rect 35909 68063 36597 68083
rect 924 68017 36611 68063
rect 924 67781 35975 68017
rect 36211 67781 36295 68017
rect 36531 67781 36611 68017
rect 924 67743 36611 67781
rect 35909 67715 36597 67743
rect 36171 67063 36859 67083
rect 452 67021 36859 67063
rect 452 66785 586 67021
rect 822 67017 36859 67021
rect 822 66785 36237 67017
rect 452 66781 36237 66785
rect 36473 66781 36557 67017
rect 36793 66781 36859 67017
rect 452 66743 36859 66781
rect 36171 66715 36859 66743
rect 36423 66063 37111 66083
rect 924 66017 37111 66063
rect 924 65781 36489 66017
rect 36725 65781 36809 66017
rect 37045 65781 37111 66017
rect 924 65743 37111 65781
rect 36423 65715 37111 65743
rect 36423 35320 37111 35345
rect 924 35279 37111 35320
rect 924 35043 36489 35279
rect 36725 35043 36809 35279
rect 37045 35043 37111 35279
rect 924 35000 37111 35043
rect 36423 34977 37111 35000
rect 36683 34320 37371 34339
rect 452 34278 37371 34320
rect 452 34042 586 34278
rect 822 34273 37371 34278
rect 822 34042 36749 34273
rect 452 34037 36749 34042
rect 36985 34037 37069 34273
rect 37305 34037 37371 34273
rect 452 34000 37371 34037
rect 36683 33971 37371 34000
rect 36936 33320 37624 33345
rect 924 33279 37624 33320
rect 924 33043 37002 33279
rect 37238 33043 37322 33279
rect 37558 33043 37624 33279
rect 924 33000 37624 33043
rect 36936 32977 37624 33000
rect 36911 2320 37599 2339
rect 924 2273 37635 2320
rect 924 2037 36977 2273
rect 37213 2037 37297 2273
rect 37533 2037 37635 2273
rect 924 2000 37635 2037
rect 36911 1971 37599 2000
rect 37195 1320 37883 1343
rect 452 1278 37883 1320
rect 452 1042 586 1278
rect 822 1277 37883 1278
rect 822 1042 37261 1277
rect 452 1041 37261 1042
rect 37497 1041 37581 1277
rect 37817 1041 37883 1277
rect 452 1000 37883 1041
rect 37195 975 37883 1000
rect 37431 320 38119 368
rect 924 302 38119 320
rect 924 66 37497 302
rect 37733 66 37817 302
rect 38053 66 38119 302
rect 924 0 38119 66
use cv3_via3_30cut  cv3_via3_30cut_0
timestamp 1563080108
transform 1 0 -566085 0 1 78451
box 566656 91154 566956 91980
use cv3_via4_2cut  cv3_via4_2cut_0
timestamp 1563080108
transform 1 0 31303 0 1 489089
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_1
timestamp 1563080108
transform 1 0 31302 0 1 470089
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_2
timestamp 1563080108
transform 1 0 31815 0 1 449090
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_3
timestamp 1563080108
transform 1 0 32327 0 1 428089
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_4
timestamp 1563080108
transform 1 0 32839 0 1 297317
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_5
timestamp 1563080108
transform 1 0 33352 0 1 264316
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_6
timestamp 1563080108
transform 1 0 33864 0 1 231341
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_7
timestamp 1563080108
transform 1 0 34375 0 1 198316
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_8
timestamp 1563080108
transform 1 0 34887 0 1 160897
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_9
timestamp 1563080108
transform 1 0 35661 0 1 99718
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_10
timestamp 1563080108
transform 1 0 36423 0 1 65715
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_11
timestamp 1563080108
transform 1 0 36423 0 1 34977
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_12
timestamp 1563080108
transform 1 0 37431 0 1 0
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_13
timestamp 1563080108
transform 1 0 37195 0 1 975
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_14
timestamp 1563080108
transform 1 0 36911 0 1 1971
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_15
timestamp 1563080108
transform 1 0 36936 0 1 32977
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_16
timestamp 1563080108
transform 1 0 36683 0 1 33971
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_17
timestamp 1563080108
transform 1 0 36171 0 1 66715
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_18
timestamp 1563080108
transform 1 0 35909 0 1 67715
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_19
timestamp 1563080108
transform 1 0 35911 0 1 98718
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_20
timestamp 1563080108
transform 1 0 35399 0 1 100716
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_21
timestamp 1563080108
transform 1 0 35147 0 1 159896
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_22
timestamp 1563080108
transform 1 0 35398 0 1 158897
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_23
timestamp 1563080108
transform 1 0 34635 0 1 197318
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_24
timestamp 1563080108
transform 1 0 34889 0 1 196317
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_25
timestamp 1563080108
transform 1 0 34123 0 1 230343
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_26
timestamp 1563080108
transform 1 0 34376 0 1 229344
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_27
timestamp 1563080108
transform 1 0 33611 0 1 263315
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_28
timestamp 1563080108
transform 1 0 33863 0 1 262317
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_29
timestamp 1563080108
transform 1 0 33099 0 1 296321
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_30
timestamp 1563080108
transform 1 0 33352 0 1 295317
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_31
timestamp 1563080108
transform 1 0 32588 0 1 427089
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_32
timestamp 1563080108
transform 1 0 32840 0 1 426091
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_33
timestamp 1563080108
transform 1 0 32075 0 1 448089
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_34
timestamp 1563080108
transform 1 0 32326 0 1 447088
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_35
timestamp 1563080108
transform 1 0 31564 0 1 469089
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_36
timestamp 1563080108
transform 1 0 31815 0 1 468089
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_37
timestamp 1563080108
transform 1 0 31051 0 1 490089
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_38
timestamp 1563080108
transform 1 0 30790 0 1 491089
box 0 0 688 368
<< properties >>
string FIXED_BBOX 0 0 38119 501877
<< end >>
