magic
tech sky130A
magscale 1 2
timestamp 1721347252
<< metal1 >>
rect 405582 59336 405782 60038
rect 405882 59336 406082 60038
rect 406182 59336 406382 60038
rect 406677 59916 407807 59944
rect 406677 59791 406725 59916
rect 406482 59616 406725 59791
rect 407761 59616 407807 59916
rect 406482 59583 407807 59616
rect 406482 59165 406682 59583
rect 422508 47562 422514 47570
rect 420993 47526 422514 47562
rect 422508 47518 422514 47526
rect 422566 47518 422572 47570
rect 420754 47158 421778 47190
rect 420754 47148 421781 47158
rect 420754 47023 420803 47148
rect 421743 47023 421781 47148
rect 420754 46988 421781 47023
rect 403880 46464 404079 46486
rect 402560 45630 402760 46056
rect 403120 45712 403156 46089
rect 403386 45797 403422 46162
rect 403663 45888 403699 46188
rect 403880 46006 403905 46464
rect 404057 46006 404079 46464
rect 403880 45980 404079 46006
rect 404186 46458 404385 46486
rect 404186 46000 404206 46458
rect 404358 46000 404385 46458
rect 420747 46173 421736 46211
rect 420747 46034 420789 46173
rect 421670 46034 421736 46173
rect 420747 46003 421736 46034
rect 404186 45980 404385 46000
rect 415700 45888 415706 45896
rect 403663 45852 415706 45888
rect 415700 45844 415706 45852
rect 415758 45888 415764 45896
rect 415758 45852 415771 45888
rect 415758 45844 415764 45852
rect 415784 45797 415790 45805
rect 403386 45761 415790 45797
rect 415784 45753 415790 45761
rect 415842 45797 415848 45805
rect 415842 45761 415857 45797
rect 415842 45753 415848 45761
rect 415868 45712 415874 45719
rect 403120 45676 415874 45712
rect 415868 45667 415874 45676
rect 415926 45712 415932 45719
rect 415926 45676 415937 45712
rect 415926 45667 415932 45676
rect 391650 45018 391672 45630
rect 392309 45018 402760 45630
rect 402906 45622 402958 45628
rect 415952 45614 415958 45621
rect 402958 45578 415958 45614
rect 402906 45564 402958 45570
rect 415952 45569 415958 45578
rect 416010 45614 416016 45621
rect 416010 45578 416018 45614
rect 416010 45569 416016 45578
rect 402908 45515 402960 45521
rect 416036 45508 416042 45514
rect 402960 45472 416042 45508
rect 402908 45457 402960 45463
rect 416036 45462 416042 45472
rect 416094 45508 416100 45514
rect 416094 45472 416102 45508
rect 416094 45462 416100 45472
rect 452721 44756 452727 44764
rect 452712 44720 452727 44756
rect 452721 44712 452727 44720
rect 452779 44756 452785 44764
rect 452779 44720 453044 44756
rect 452779 44712 452785 44720
rect 446714 44672 446720 44680
rect 446698 44636 446720 44672
rect 446714 44628 446720 44636
rect 446772 44672 446778 44680
rect 446772 44636 453044 44672
rect 446772 44628 446778 44636
rect 452559 44588 452565 44596
rect 452550 44552 452565 44588
rect 452559 44544 452565 44552
rect 452617 44588 452623 44596
rect 452617 44552 453044 44588
rect 452617 44544 452623 44552
rect 446878 44504 446884 44512
rect 446862 44468 446884 44504
rect 446878 44460 446884 44468
rect 446936 44504 446942 44512
rect 446936 44468 453044 44504
rect 446936 44460 446942 44468
rect 452399 44420 452405 44428
rect 452392 44384 452405 44420
rect 452399 44376 452405 44384
rect 452457 44420 452463 44428
rect 452457 44384 453044 44420
rect 452457 44376 452463 44384
rect 447037 44336 447043 44344
rect 447019 44300 447043 44336
rect 447037 44292 447043 44300
rect 447095 44336 447101 44344
rect 447095 44300 453044 44336
rect 447095 44292 447101 44300
rect 452237 44252 452243 44260
rect 452235 44216 452243 44252
rect 452237 44208 452243 44216
rect 452295 44252 452301 44260
rect 452295 44216 453044 44252
rect 452295 44208 452301 44216
rect 447201 44168 447207 44176
rect 447177 44132 447207 44168
rect 447201 44124 447207 44132
rect 447259 44168 447265 44176
rect 447259 44132 453044 44168
rect 447259 44124 447265 44132
rect 452082 44084 452088 44092
rect 452080 44048 452088 44084
rect 452082 44040 452088 44048
rect 452140 44084 452146 44092
rect 452140 44048 453044 44084
rect 452140 44040 452146 44048
rect 447354 44000 447365 44008
rect 447345 43964 447365 44000
rect 447354 43956 447365 43964
rect 447417 44000 447423 44008
rect 447417 43964 453044 44000
rect 447417 43956 447423 43964
rect 451914 43872 451920 43924
rect 451972 43916 451978 43924
rect 451972 43880 453044 43916
rect 451972 43872 451978 43880
rect 447518 43832 447524 43840
rect 447507 43796 447524 43832
rect 447518 43788 447524 43796
rect 447576 43832 447582 43840
rect 447576 43796 453044 43832
rect 447576 43788 447582 43796
rect 451759 43748 451765 43756
rect 451754 43712 451765 43748
rect 451759 43704 451765 43712
rect 451817 43748 451823 43756
rect 451817 43712 453044 43748
rect 451817 43704 451823 43712
rect 447682 43664 447688 43672
rect 447664 43628 447688 43664
rect 447682 43620 447688 43628
rect 447740 43664 447746 43672
rect 447740 43628 453044 43664
rect 447740 43620 447746 43628
rect 451597 43580 451603 43588
rect 451590 43544 451603 43580
rect 451597 43536 451603 43544
rect 451655 43580 451661 43588
rect 451655 43544 453044 43580
rect 451655 43536 451661 43544
rect 447840 43496 447846 43504
rect 447819 43460 447846 43496
rect 447840 43452 447846 43460
rect 447898 43496 447904 43504
rect 447898 43460 453044 43496
rect 447898 43452 447904 43460
rect 457038 30024 457238 30030
rect 457038 28017 457238 29824
rect 458027 30010 458227 30016
rect 458027 28017 458227 29810
rect 458462 28016 458538 28967
rect 458753 28002 458829 28953
<< via1 >>
rect 406725 59616 407761 59916
rect 422514 47518 422566 47570
rect 420803 47023 421743 47148
rect 403905 46006 404057 46464
rect 404206 46000 404358 46458
rect 420789 46034 421670 46173
rect 415706 45844 415758 45896
rect 415790 45753 415842 45805
rect 415874 45667 415926 45719
rect 391672 45018 392309 45630
rect 402906 45570 402958 45622
rect 415958 45569 416010 45621
rect 402908 45463 402960 45515
rect 416042 45462 416094 45514
rect 452727 44712 452779 44764
rect 446720 44628 446772 44680
rect 452565 44544 452617 44596
rect 446884 44460 446936 44512
rect 452405 44376 452457 44428
rect 447043 44292 447095 44344
rect 452243 44208 452295 44260
rect 447207 44124 447259 44176
rect 452088 44040 452140 44092
rect 447365 43956 447417 44008
rect 451920 43872 451972 43924
rect 447524 43788 447576 43840
rect 451765 43704 451817 43756
rect 447688 43620 447740 43672
rect 451603 43536 451655 43588
rect 447846 43452 447898 43504
rect 457038 29824 457238 30024
rect 458027 29810 458227 30010
<< metal2 >>
rect 405578 60978 405749 60987
rect 405578 60398 405749 60807
rect 405907 60610 406050 66606
rect 406227 60550 406370 66546
rect 422027 60976 422210 60985
rect 406677 59916 407807 59944
rect 406677 59616 406725 59916
rect 407761 59616 407807 59916
rect 406677 59583 407807 59616
rect 387066 54146 387138 54316
rect 387080 49530 387116 54146
rect 391304 53896 391358 54104
rect 385998 49494 387116 49530
rect 385998 44160 386034 49494
rect 385998 44124 386234 44160
rect 385241 43716 386119 43750
rect 385241 43242 385274 43716
rect 386087 43242 386119 43716
rect 385241 43211 386119 43242
rect 386198 42399 386234 44124
rect 385408 42363 386234 42399
rect 384012 41614 385956 41662
rect 384012 41169 384078 41614
rect 385891 41169 385956 41614
rect 384012 41112 385956 41169
rect 367620 40310 368082 40315
rect 367616 40203 367625 40310
rect 367732 40203 368082 40310
rect 391314 40264 391350 53896
rect 385529 40228 391350 40264
rect 391672 45630 392309 45646
rect 401933 45507 401969 46594
rect 402220 45614 402256 46470
rect 403880 46464 404079 46486
rect 403880 46006 403905 46464
rect 404057 46006 404079 46464
rect 403880 45980 404079 46006
rect 404186 46458 404385 46486
rect 404186 46000 404206 46458
rect 404358 46000 404385 46458
rect 404186 45980 404385 46000
rect 415714 45902 415750 60574
rect 415706 45896 415758 45902
rect 415706 45838 415758 45844
rect 415714 45834 415750 45838
rect 415798 45811 415834 60574
rect 415790 45805 415842 45811
rect 415790 45747 415842 45753
rect 415798 45741 415834 45747
rect 415882 45725 415918 60574
rect 415874 45719 415926 45725
rect 415874 45661 415926 45667
rect 415882 45652 415918 45661
rect 415966 45627 416002 60574
rect 402900 45614 402906 45622
rect 402220 45578 402906 45614
rect 402900 45570 402906 45578
rect 402958 45570 402964 45622
rect 415958 45621 416010 45627
rect 415958 45563 416010 45569
rect 415966 45558 416002 45563
rect 416050 45520 416086 60574
rect 421035 51919 421805 51943
rect 421035 51916 421070 51919
rect 420956 51773 421070 51916
rect 421767 51773 421805 51919
rect 420956 51748 421805 51773
rect 421035 51738 421805 51748
rect 422027 51471 422210 60793
rect 422492 59522 422580 59788
rect 420904 51288 422210 51471
rect 416981 49325 417583 49462
rect 402902 45507 402908 45515
rect 401933 45471 402908 45507
rect 402902 45463 402908 45471
rect 402960 45463 402966 45515
rect 416042 45514 416094 45520
rect 416042 45456 416094 45462
rect 416050 45451 416086 45456
rect 367620 40198 368082 40203
rect 391672 39723 392309 45018
rect 385452 39086 392309 39723
rect 392687 29414 392827 44520
rect 416981 44430 417118 49325
rect 421021 48814 422062 48919
rect 420994 48487 421764 48507
rect 420994 48341 421046 48487
rect 421743 48341 421764 48487
rect 420994 48317 421764 48341
rect 420754 47158 421778 47190
rect 420754 47148 421781 47158
rect 420754 47023 420803 47148
rect 421743 47023 421781 47148
rect 420754 46988 421781 47023
rect 420747 46173 421736 46211
rect 420747 46034 420789 46173
rect 421670 46034 421736 46173
rect 420747 46003 421736 46034
rect 421950 44616 422062 48814
rect 422522 47576 422558 59522
rect 422514 47570 422566 47576
rect 422514 47512 422566 47518
rect 430508 37750 430580 60082
rect 430094 37678 430580 37750
rect 430608 36998 430676 60082
rect 430084 36930 430676 36998
rect 393739 32731 395092 32753
rect 393739 32474 393779 32731
rect 394848 32474 395092 32731
rect 430724 32645 430760 60082
rect 430265 32609 430760 32645
rect 393739 32443 395092 32474
rect 430255 31890 430749 31916
rect 430715 31573 430749 31890
rect 430255 31541 430749 31573
rect 430808 31114 430844 60082
rect 446720 45172 446789 45187
rect 436476 44757 436556 45046
rect 446720 44680 446789 44838
rect 446772 44628 446789 44680
rect 446720 44619 446789 44628
rect 446880 45172 446949 45187
rect 446880 44512 446949 44838
rect 446880 44460 446884 44512
rect 446936 44460 446949 44512
rect 446880 44453 446949 44460
rect 447040 45172 447109 45187
rect 447040 44344 447109 44838
rect 447040 44292 447043 44344
rect 447095 44292 447109 44344
rect 447040 44273 447109 44292
rect 447200 45172 447269 45187
rect 447200 44176 447269 44838
rect 447200 44124 447207 44176
rect 447259 44124 447269 44176
rect 447200 44113 447269 44124
rect 447360 45172 447429 45187
rect 447360 44008 447429 44838
rect 447360 43956 447365 44008
rect 447417 43956 447429 44008
rect 447360 43949 447429 43956
rect 447520 45172 447589 45187
rect 447520 43840 447589 44838
rect 447520 43788 447524 43840
rect 447576 43788 447589 43840
rect 447520 43774 447589 43788
rect 447680 45172 447749 45187
rect 447680 43672 447749 44838
rect 447680 43620 447688 43672
rect 447740 43620 447749 43672
rect 447680 43607 447749 43620
rect 447840 45172 447909 45187
rect 447840 43504 447909 44838
rect 451596 45175 451665 45190
rect 451596 43588 451665 44841
rect 451756 45175 451825 45190
rect 451756 43756 451825 44841
rect 451916 45175 451985 45190
rect 451916 43924 451985 44841
rect 452076 45175 452145 45190
rect 452076 44092 452145 44841
rect 452236 45175 452305 45190
rect 452236 44260 452305 44841
rect 452396 45175 452465 45190
rect 452396 44428 452465 44841
rect 452556 45175 452625 45190
rect 452556 44596 452625 44841
rect 452716 45175 452785 45190
rect 452716 44764 452785 44841
rect 452716 44712 452727 44764
rect 452779 44712 452785 44764
rect 452716 44697 452785 44712
rect 452556 44544 452565 44596
rect 452617 44544 452625 44596
rect 452556 44532 452625 44544
rect 452396 44376 452405 44428
rect 452457 44376 452465 44428
rect 452396 44366 452465 44376
rect 452236 44208 452243 44260
rect 452295 44208 452305 44260
rect 452236 44190 452305 44208
rect 452076 44040 452088 44092
rect 452140 44040 452145 44092
rect 452076 44028 452145 44040
rect 451916 43872 451920 43924
rect 451972 43872 451985 43924
rect 451916 43864 451985 43872
rect 451756 43704 451765 43756
rect 451817 43704 451825 43756
rect 451756 43691 451825 43704
rect 451596 43536 451603 43588
rect 451655 43536 451665 43588
rect 451596 43519 451665 43536
rect 447840 43452 447846 43504
rect 447898 43452 447909 43504
rect 447840 43439 447909 43452
rect 430214 31078 430844 31114
rect 457038 31225 457238 31234
rect 457038 30024 457238 31025
rect 458027 30778 458227 30787
rect 457032 29824 457038 30024
rect 457238 29824 457244 30024
rect 458027 30010 458227 30578
rect 458021 29810 458027 30010
rect 458227 29810 458233 30010
rect 459366 29925 459566 29934
rect 392687 29318 394379 29414
rect 392020 29084 394378 29116
rect 392020 28615 392065 29084
rect 392969 28615 394378 29084
rect 392020 28577 394378 28615
rect 459366 27994 459566 29725
rect 464230 29833 464430 29842
rect 464230 27994 464430 29633
rect 459688 22181 460660 23289
rect 459688 21958 459730 22181
rect 460617 21958 460660 22181
rect 459688 21920 460660 21958
rect 463140 22162 464113 23289
rect 463140 21939 463174 22162
rect 464061 21939 464113 22162
rect 463140 21920 464113 21939
<< via2 >>
rect 405578 60807 405749 60978
rect 422027 60793 422210 60976
rect 406725 59616 407761 59916
rect 385274 43242 386087 43716
rect 384078 41169 385891 41614
rect 367625 40203 367732 40310
rect 403905 46006 404057 46464
rect 404206 46000 404358 46458
rect 421070 51773 421767 51919
rect 421046 48341 421743 48487
rect 420803 47023 421743 47148
rect 420789 46034 421670 46173
rect 393779 32474 394848 32731
rect 430108 31573 430715 31890
rect 446720 44838 446789 45172
rect 446880 44838 446949 45172
rect 447040 44838 447109 45172
rect 447200 44838 447269 45172
rect 447360 44838 447429 45172
rect 447520 44838 447589 45172
rect 447680 44838 447749 45172
rect 447840 44838 447909 45172
rect 451596 44841 451665 45175
rect 451756 44841 451825 45175
rect 451916 44841 451985 45175
rect 452076 44841 452145 45175
rect 452236 44841 452305 45175
rect 452396 44841 452465 45175
rect 452556 44841 452625 45175
rect 452716 44841 452785 45175
rect 457038 31025 457238 31225
rect 458027 30578 458227 30778
rect 459366 29725 459566 29925
rect 392065 28615 392969 29084
rect 464230 29633 464430 29833
rect 459730 21958 460617 22181
rect 463174 21939 464061 22162
<< metal3 >>
rect 405573 60978 405754 60983
rect 422022 60978 422215 60981
rect 405573 60807 405578 60978
rect 405749 60976 422228 60978
rect 405749 60807 422027 60976
rect 405573 60802 405754 60807
rect 413700 60760 415496 60807
rect 422022 60793 422027 60807
rect 422210 60807 422228 60976
rect 422210 60793 422215 60807
rect 422022 60788 422215 60793
rect 413700 60480 413748 60760
rect 415458 60480 415496 60760
rect 413700 60440 415496 60480
rect 405417 59916 406546 59943
rect 406677 59916 407807 59944
rect 405417 59616 405465 59916
rect 406501 59616 406725 59916
rect 407761 59616 407807 59916
rect 405417 59583 406546 59616
rect 406677 59583 407807 59616
rect 421035 51919 421805 51943
rect 421035 51773 421070 51919
rect 421767 51773 421805 51919
rect 421035 51738 421805 51773
rect 421004 48487 421774 48515
rect 421004 48341 421046 48487
rect 421743 48341 421774 48487
rect 421004 48310 421774 48341
rect 420754 47158 421778 47190
rect 420754 47148 421781 47158
rect 420754 47023 420803 47148
rect 421743 47023 421781 47148
rect 420754 46988 421781 47023
rect 403880 46464 404079 46486
rect 403880 46006 403905 46464
rect 404057 46006 404079 46464
rect 403880 45978 404079 46006
rect 404186 46458 404385 46486
rect 404186 46000 404206 46458
rect 404358 46000 404385 46458
rect 420747 46173 421736 46211
rect 420747 46034 420789 46173
rect 421670 46034 421736 46173
rect 420747 46003 421736 46034
rect 403756 45940 404086 45978
rect 402878 45342 403415 45397
rect 402878 44613 402922 45342
rect 403374 44767 403415 45342
rect 403756 44919 403806 45940
rect 404042 44919 404086 45940
rect 403756 44879 404086 44919
rect 403880 44875 404079 44879
rect 404186 44767 404385 46000
rect 446715 45172 446795 45218
rect 446715 44838 446720 45172
rect 446789 44838 446795 45172
rect 446715 44832 446795 44838
rect 446875 45172 446955 45218
rect 446875 44838 446880 45172
rect 446949 44838 446955 45172
rect 446875 44832 446955 44838
rect 447035 45172 447115 45218
rect 447035 44838 447040 45172
rect 447109 44838 447115 45172
rect 447035 44832 447115 44838
rect 447195 45172 447275 45218
rect 447195 44838 447200 45172
rect 447269 44838 447275 45172
rect 447195 44832 447275 44838
rect 447355 45172 447435 45218
rect 447355 44838 447360 45172
rect 447429 44838 447435 45172
rect 447355 44832 447435 44838
rect 447515 45172 447595 45218
rect 447515 44838 447520 45172
rect 447589 44838 447595 45172
rect 447515 44832 447595 44838
rect 447675 45172 447755 45218
rect 447675 44838 447680 45172
rect 447749 44838 447755 45172
rect 447675 44832 447755 44838
rect 447835 45172 447915 45218
rect 447835 44838 447840 45172
rect 447909 44838 447915 45172
rect 447835 44832 447915 44838
rect 451591 45175 451671 45192
rect 451591 44841 451596 45175
rect 451665 44841 451671 45175
rect 451591 44835 451671 44841
rect 451751 45175 451831 45192
rect 451751 44841 451756 45175
rect 451825 44841 451831 45175
rect 451751 44835 451831 44841
rect 451911 45175 451991 45192
rect 451911 44841 451916 45175
rect 451985 44841 451991 45175
rect 451911 44835 451991 44841
rect 452071 45175 452151 45192
rect 452071 44841 452076 45175
rect 452145 44841 452151 45175
rect 452071 44835 452151 44841
rect 452231 45175 452311 45192
rect 452231 44841 452236 45175
rect 452305 44841 452311 45175
rect 452231 44835 452311 44841
rect 452391 45175 452471 45192
rect 452391 44841 452396 45175
rect 452465 44841 452471 45175
rect 452391 44835 452471 44841
rect 452551 45175 452631 45192
rect 452551 44841 452556 45175
rect 452625 44841 452631 45175
rect 452551 44835 452631 44841
rect 452711 44841 452716 44966
rect 452785 44841 452791 44966
rect 452711 44835 452791 44841
rect 403374 44613 404385 44767
rect 421907 44652 436556 44757
rect 402878 44569 404385 44613
rect 402886 44568 404385 44569
rect 367620 44430 390179 44547
rect 367620 40310 367737 44430
rect 390062 44401 390179 44430
rect 444172 44401 444956 44496
rect 390062 44284 455685 44401
rect 455802 44284 455808 44401
rect 444172 44224 444956 44284
rect 385241 43716 386119 43750
rect 385241 43242 385274 43716
rect 386087 43242 386119 43716
rect 385241 43211 386119 43242
rect 384012 41614 385956 41662
rect 384012 41169 384078 41614
rect 385891 41169 385956 41614
rect 384012 41112 385956 41169
rect 367620 40203 367625 40310
rect 367732 40203 367737 40310
rect 367620 40198 367737 40203
rect 389683 32738 394881 32754
rect 389683 32467 389701 32738
rect 391045 32731 394881 32738
rect 391045 32474 393779 32731
rect 394848 32474 394881 32731
rect 391045 32467 394881 32474
rect 389683 32447 394881 32467
rect 430070 31895 433193 31918
rect 430070 31890 432505 31895
rect 430070 31573 430108 31890
rect 430715 31573 432505 31890
rect 430070 31571 432505 31573
rect 433161 31571 433193 31895
rect 430070 31545 433193 31571
rect 457033 31225 457243 31230
rect 457033 31025 457038 31225
rect 457238 31025 461411 31225
rect 461611 31025 461617 31225
rect 457033 31020 457243 31025
rect 458022 30778 458232 30783
rect 458022 30578 458027 30778
rect 458227 30578 460722 30778
rect 460922 30578 460928 30778
rect 458022 30573 458232 30578
rect 459361 29925 459571 29930
rect 459361 29725 459366 29925
rect 459566 29725 462159 29925
rect 462359 29725 462365 29925
rect 464225 29833 464435 29838
rect 459361 29720 459571 29725
rect 462908 29633 462914 29833
rect 463114 29633 464230 29833
rect 464430 29633 464435 29833
rect 464225 29628 464435 29633
rect 391405 29084 393015 29129
rect 391405 28593 391451 29084
rect 392975 28593 393015 29084
rect 391405 28550 393015 28593
rect 459688 22193 460667 22218
rect 458965 22181 460667 22193
rect 458965 22158 459730 22181
rect 455685 22157 459730 22158
rect 455680 22042 455686 22157
rect 455801 22042 459730 22157
rect 455685 22041 459730 22042
rect 458965 21999 459730 22041
rect 459688 21958 459730 21999
rect 460617 21958 460667 22181
rect 459688 21920 460667 21958
rect 463140 22162 464099 22186
rect 463140 21939 463174 22162
rect 464061 22147 464099 22162
rect 464061 21953 464825 22147
rect 464061 21939 464099 21953
rect 463140 21920 464099 21939
<< via3 >>
rect 413748 60480 415458 60760
rect 405465 59616 406501 59916
rect 421070 51773 421767 51919
rect 421046 48341 421743 48487
rect 420803 47023 421743 47148
rect 420789 46034 421670 46173
rect 402922 44613 403374 45342
rect 403806 44919 404042 45940
rect 455685 44284 455802 44401
rect 385274 43242 386087 43716
rect 384078 41169 385891 41614
rect 389701 32467 391045 32738
rect 432505 31571 433161 31895
rect 461411 31025 461611 31225
rect 460722 30578 460922 30778
rect 462159 29725 462359 29925
rect 462914 29633 463114 29833
rect 391451 28615 392065 29084
rect 392065 28615 392969 29084
rect 392969 28615 392975 29084
rect 391451 28593 392975 28615
rect 455686 22042 455801 22157
<< metal4 >>
rect 385422 70030 386100 70143
rect 385422 68868 385480 70030
rect 386034 68868 386100 70030
rect 384357 67952 385102 68058
rect 384357 66822 384412 67952
rect 385024 66822 385102 67952
rect 382912 53463 383955 53537
rect 382912 50614 382998 53463
rect 383893 50614 383955 53463
rect 382912 50530 383955 50614
rect 368182 45515 369817 45667
rect 368182 45451 368294 45515
rect 368180 44750 368294 45451
rect 369665 44750 369817 45515
rect 368180 44591 369817 44750
rect 368180 43841 368577 44591
rect 383168 39215 383713 50530
rect 384357 41662 385102 66822
rect 385422 43750 386100 68868
rect 404527 70054 405080 70078
rect 404527 68864 404568 70054
rect 405032 68864 405080 70054
rect 399435 67992 399974 68095
rect 399435 66802 399468 67992
rect 399932 66802 399974 67992
rect 385241 43716 386100 43750
rect 385241 43242 385274 43716
rect 386087 43242 386100 43716
rect 385241 43211 386100 43242
rect 389684 53468 391062 53564
rect 389684 50582 389744 53468
rect 390995 50582 391062 53468
rect 399435 53451 399974 66802
rect 404527 53483 405080 68864
rect 429864 70050 430192 70121
rect 429864 68838 429882 70050
rect 430167 68838 430192 70050
rect 422531 65770 423281 65881
rect 422531 63924 422572 65770
rect 423220 63924 423281 65770
rect 421472 63012 422241 63052
rect 421472 61166 421520 63012
rect 422168 61166 422241 63012
rect 413700 60760 415496 60810
rect 413700 60480 413748 60760
rect 415458 60480 415496 60760
rect 413700 60440 415496 60480
rect 421472 60080 422241 61166
rect 422531 60769 423281 63924
rect 422531 60082 429638 60769
rect 405417 59916 406547 59944
rect 405417 59616 405465 59916
rect 406501 59616 406547 59916
rect 405417 59583 406547 59616
rect 399435 52912 403417 53451
rect 384012 41614 385956 41662
rect 384012 41169 384078 41614
rect 385891 41169 385956 41614
rect 384012 41112 385956 41169
rect 372113 38670 383713 39215
rect 389684 32738 391062 50582
rect 389684 32467 389701 32738
rect 391045 32467 391062 32738
rect 389684 32431 391062 32467
rect 391399 48413 392808 48502
rect 391399 45614 391494 48413
rect 392733 45614 392808 48413
rect 391399 29129 392808 45614
rect 402878 45342 403417 52912
rect 402878 44613 402922 45342
rect 403374 44613 403417 45342
rect 403760 52930 405080 53483
rect 403760 45940 404313 52930
rect 403760 44919 403806 45940
rect 404042 44919 404313 45940
rect 405446 48473 406518 59583
rect 414900 59311 422241 60080
rect 422518 60014 429638 60082
rect 414900 52381 415669 59311
rect 414900 51919 422027 52381
rect 414900 51773 421070 51919
rect 421767 51773 422027 51919
rect 414900 51612 422027 51773
rect 428888 50307 429638 60014
rect 421022 49557 429638 50307
rect 421022 48515 421772 49557
rect 405446 45583 405504 48473
rect 406457 45583 406518 48473
rect 421004 48487 421774 48515
rect 421004 48341 421046 48487
rect 421743 48341 421774 48487
rect 421004 48310 421774 48341
rect 429864 47261 430192 68838
rect 477949 70010 478802 70070
rect 477949 68878 478016 70010
rect 478718 68878 478802 70010
rect 420743 47148 430192 47261
rect 420743 47023 420803 47148
rect 421743 47023 430192 47148
rect 420743 46933 430192 47023
rect 430337 67982 430665 68016
rect 430337 66778 430355 67982
rect 430640 66778 430665 67982
rect 430337 46281 430665 66778
rect 476762 67968 477619 68060
rect 476762 66836 476844 67968
rect 477546 66836 477619 67968
rect 476762 59794 477619 66836
rect 473864 58834 477619 59794
rect 477949 59826 478802 68878
rect 484412 70065 484854 70217
rect 484412 68863 484446 70065
rect 484801 68863 484854 70065
rect 477949 58866 481361 59826
rect 477949 58865 478013 58866
rect 420728 46173 430665 46281
rect 420728 46034 420789 46173
rect 421670 46034 430665 46173
rect 420728 45953 430665 46034
rect 480401 45966 481361 58866
rect 405446 45522 406518 45583
rect 403760 44879 404313 44919
rect 402878 44550 403417 44613
rect 393134 29721 393549 38162
rect 432479 31895 433187 45918
rect 474624 45006 481361 45966
rect 455684 44401 455803 44402
rect 455684 44284 455685 44401
rect 455802 44284 455803 44401
rect 455684 44283 455803 44284
rect 432479 31571 432505 31895
rect 433161 31571 433187 31895
rect 432479 31545 433187 31571
rect 391399 29084 393015 29129
rect 391399 28593 391451 29084
rect 392975 28593 393015 29084
rect 391399 28566 393015 28593
rect 391405 28550 393015 28566
rect 393221 25358 393548 29721
rect 455685 22157 455802 44283
rect 484412 43935 484854 68863
rect 460597 43493 484854 43935
rect 485114 67986 485556 68245
rect 485114 66784 485146 67986
rect 485501 66784 485556 67986
rect 460597 30778 461039 43493
rect 485114 43233 485556 66784
rect 460597 30578 460722 30778
rect 460922 30578 461039 30778
rect 460597 23087 461039 30578
rect 461299 42791 485556 43233
rect 485860 65778 486302 65947
rect 485860 63913 485890 65778
rect 486259 63913 486302 65778
rect 461299 31225 461741 42791
rect 485860 42487 486302 63913
rect 461299 31025 461411 31225
rect 461611 31025 461741 31225
rect 461299 23189 461741 31025
rect 462045 42045 486302 42487
rect 486623 63001 487065 63242
rect 486623 61149 486664 63001
rect 487021 61149 487065 63001
rect 462045 29925 462487 42045
rect 486623 41724 487065 61149
rect 462045 29725 462159 29925
rect 462359 29725 462487 29925
rect 462045 23204 462487 29725
rect 462808 41282 487065 41724
rect 462808 29833 463250 41282
rect 462808 29633 462914 29833
rect 463114 29633 463250 29833
rect 462808 23135 463250 29633
rect 455685 22042 455686 22157
rect 455801 22042 455802 22157
rect 455685 22041 455802 22042
<< via4 >>
rect 385480 68868 386034 70030
rect 384412 66822 385024 67952
rect 382998 50614 383893 53463
rect 368294 44750 369665 45515
rect 404568 68864 405032 70054
rect 399468 66802 399932 67992
rect 389744 50582 390995 53468
rect 429882 68838 430167 70050
rect 422572 63924 423220 65770
rect 421520 61166 422168 63012
rect 413748 60480 415458 60760
rect 391494 45614 392733 48413
rect 405504 45583 406457 48473
rect 478016 68878 478718 70010
rect 430355 66778 430640 67982
rect 476844 66836 477546 67968
rect 484446 68863 484801 70065
rect 485146 66784 485501 67986
rect 485890 63913 486259 65778
rect 486664 61149 487021 63001
<< metal5 >>
rect 367122 70065 487354 70090
rect 367122 70054 484446 70065
rect 367122 70030 404568 70054
rect 367122 68868 385480 70030
rect 386034 68868 404568 70030
rect 367122 68864 404568 68868
rect 405032 70050 484446 70054
rect 405032 68864 429882 70050
rect 367122 68838 429882 68864
rect 430167 70010 484446 70050
rect 430167 68878 478016 70010
rect 478718 68878 484446 70010
rect 430167 68863 484446 68878
rect 484801 68863 487354 70065
rect 430167 68838 487354 68863
rect 367122 68814 487354 68838
rect 367076 67992 487354 68024
rect 367076 67952 399468 67992
rect 367076 66822 384412 67952
rect 385024 66822 399468 67952
rect 367076 66802 399468 66822
rect 399932 67986 487354 67992
rect 399932 67982 485146 67986
rect 399932 66802 430355 67982
rect 367076 66778 430355 66802
rect 430640 67968 485146 67982
rect 430640 66836 476844 67968
rect 477546 66836 485146 67968
rect 430640 66784 485146 66836
rect 485501 66784 487354 67986
rect 430640 66778 487354 66784
rect 367076 66748 487354 66778
rect 367050 65778 487354 65820
rect 367050 65770 485890 65778
rect 367050 63924 422572 65770
rect 423220 63924 485890 65770
rect 367050 63913 485890 63924
rect 486259 63913 487354 65778
rect 367050 63878 487354 63913
rect 367098 63012 487354 63054
rect 367098 61166 421520 63012
rect 422168 63001 487354 63012
rect 422168 61166 486664 63001
rect 367098 61149 486664 61166
rect 487021 61149 487354 63001
rect 367098 61112 487354 61149
rect 413700 60760 415496 60786
rect 413700 60480 413748 60760
rect 415458 60480 415496 60760
rect 413700 60440 415496 60480
rect 415095 57822 415495 60440
rect 415095 57384 427817 57822
rect 415095 54589 415495 57384
rect 429227 56295 430088 56297
rect 415939 55885 430088 56295
rect 415095 54151 427764 54589
rect 366986 53468 391206 53534
rect 366986 53463 389744 53468
rect 366986 50614 382998 53463
rect 383893 50614 389744 53463
rect 366986 50582 389744 50614
rect 390995 50582 391206 53468
rect 429227 53031 430088 55885
rect 415939 52621 430088 53031
rect 366986 50534 391206 50582
rect 429227 48534 430088 52621
rect 366986 48473 487354 48534
rect 366986 48413 405504 48473
rect 366986 45614 391494 48413
rect 392733 45614 405504 48413
rect 366986 45583 405504 45614
rect 406457 45583 487354 48473
rect 366986 45534 487354 45583
rect 368182 45515 369817 45534
rect 368182 44750 368294 45515
rect 369665 44750 369817 45515
rect 368182 44591 369817 44750
use cv3_via2_36cut  cv3_via2_36cut_222
timestamp 1719173892
transform 1 0 -133419 0 1 -47639
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_223
timestamp 1719173892
transform 1 0 -162625 0 1 -48017
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_224
timestamp 1719173892
transform 1 0 -139036 0 1 -48028
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_225
timestamp 1719173892
transform 1 0 -119549 0 1 -47621
box 555256 92202 556228 92502
use cv3_via_30cut  cv3_via_30cut_12
timestamp 1719247715
transform 1 0 391188 0 1 -44926
box 14334 104924 14594 105610
use cv3_via_30cut  cv3_via_30cut_13
timestamp 1719247715
transform 1 0 391849 0 1 -44917
box 14334 104924 14594 105610
use cv3_via_30cut  cv3_via_30cut_14
timestamp 1719247715
transform 1 0 391520 0 1 -44919
box 14334 104924 14594 105610
use isolated_switch_xlarge  isolated_switch_xlarge_0 ../ip/sky130_ef_ip__analog_switches/mag
timestamp 1719257891
transform 0 -1 458356 -1 0 28707
box 660 -6310 5486 1338
use simple_analog_mux_sel1v8  simple_analog_mux_sel1v8_1 ../ip/sky130_ef_ip__analog_switches/mag
timestamp 1719277428
transform -1 0 421022 0 -1 49627
box -46 -2540 3538 3648
use sky130_ak_ip__cmos_vref  sky130_ak_ip__cmos_vref_0 ../ip/sky130_ak_ip__cmos_vref/mag
timestamp 1721067183
transform 0 -1 395482 1 0 37455
box 8587 -19903 21921 206
use sky130_am_ip__ldo_01v8  sky130_am_ip__ldo_01v8_0 ../ip/sky130_am_ip__ldo_01v8/mag
timestamp 1721052427
transform 0 1 378665 -1 0 48529
box 4253 -10775 28439 6899
use sky130_cw_ip__bandgap  sky130_cw_ip__bandgap_0 ../ip/sky130_cw_ip/mag
timestamp 1715625863
transform -1 0 474518 0 1 44954
box -5734 12 42048 14837
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_1
array 0 1 3268 0 4 2588
timestamp 1721093827
transform 0 1 417124 -1 0 57339
box -1349 -1081 1371 1081
use sky130_sw_ip__bgrref_por  sky130_sw_ip__bgrref_por_0 ../ip/sky130_sw_ip__bgrref_por/mag
timestamp 1721154165
transform 1 0 390789 0 1 321922
box 2359 -300396 39662 -277894
<< labels >>
flabel metal5 367470 46090 370116 48014 0 FreeSans 4800 0 0 0 vssio
port 1 nsew
flabel metal5 367390 51088 370170 53332 0 FreeSans 4800 0 0 0 vddio
port 0 nsew
flabel metal5 367230 66874 369822 67890 0 FreeSans 3200 0 0 0 vssd0
port 2 nsew
flabel metal5 367256 69000 369848 70016 0 FreeSans 3200 0 0 0 vccd0
port 3 nsew
flabel metal5 367342 64120 369672 65674 0 FreeSans 4800 0 0 0 vdda0
port 4 nsew
flabel metal5 367294 61354 369624 62908 0 FreeSans 4800 0 0 0 vssa0
port 5 nsew
flabel metal2 391304 53896 391358 54104 0 FreeSans 320 90 0 0 ldo_ref_sel
port 6 nsew
flabel metal2 387066 54146 387138 54316 0 FreeSans 320 90 0 0 ldo_ena
port 7 nsew
flabel metal3 444172 44224 444956 44496 0 FreeSans 800 0 0 0 vbg
port 8 nsew
flabel metal1 452779 44720 453044 44756 0 FreeSans 320 0 0 0 bandgap_trim[0]
port 9 nsew
flabel metal1 452744 44636 453044 44672 0 FreeSans 320 0 0 0 bandgap_trim[1]
port 10 nsew
flabel metal1 452744 44552 453044 44588 0 FreeSans 320 0 0 0 bandgap_trim[2]
port 11 nsew
flabel metal1 452744 44468 453044 44504 0 FreeSans 320 0 0 0 bandgap_trim[3]
port 12 nsew
flabel metal1 452744 44384 453044 44420 0 FreeSans 320 0 0 0 bandgap_trim[4]
port 13 nsew
flabel metal1 452744 44300 453044 44336 0 FreeSans 320 0 0 0 bandgap_trim[5]
port 14 nsew
flabel metal1 452744 44216 453044 44252 0 FreeSans 320 0 0 0 bandgap_trim[6]
port 15 nsew
flabel metal1 452744 44132 453044 44168 0 FreeSans 320 0 0 0 bandgap_trim[7]
port 16 nsew
flabel metal1 452744 44048 453044 44084 0 FreeSans 320 0 0 0 bandgap_trim[8]
port 17 nsew
flabel metal1 452744 43964 453044 44000 0 FreeSans 320 0 0 0 bandgap_trim[9]
port 18 nsew
flabel metal1 452744 43880 453044 43916 0 FreeSans 320 0 0 0 bandgap_trim[10]
port 19 nsew
flabel metal1 452744 43796 453044 43832 0 FreeSans 320 0 0 0 bandgap_trim[11]
port 20 nsew
flabel metal1 452744 43712 453044 43748 0 FreeSans 320 0 0 0 bandgap_trim[12]
port 21 nsew
flabel metal1 452744 43628 453044 43664 0 FreeSans 320 0 0 0 bandgap_trim[13]
port 22 nsew
flabel metal1 452744 43544 453044 43580 0 FreeSans 320 0 0 0 bandgap_trim[14]
port 23 nsew
flabel metal1 452744 43460 453044 43496 0 FreeSans 320 0 0 0 bandgap_trim[15]
port 24 nsew
flabel metal2 422492 59522 422580 59788 0 FreeSans 320 90 0 0 bandgap_sel
port 25 nsew
flabel metal2 430508 59782 430580 60082 0 FreeSans 320 90 0 0 porb_h[0]
port 26 nsew
flabel metal2 430608 59782 430676 60082 0 FreeSans 320 90 0 0 porb_h[1]
port 27 nsew
flabel metal2 430724 59782 430760 60082 0 FreeSans 320 90 0 0 porb
port 28 nsew
flabel metal2 430808 59782 430844 60082 0 FreeSans 320 90 0 0 por
port 29 nsew
flabel metal2 415714 60274 415750 60574 0 FreeSans 320 90 0 0 bandgap_ena
port 30 nsew
flabel metal2 415798 60274 415834 60574 0 FreeSans 320 90 0 0 bandgap_trim[3]
port 32 nsew
flabel metal2 415882 60274 415918 60574 0 FreeSans 320 90 0 0 bandgap_trim[2]
port 33 nsew
flabel metal2 415966 60274 416002 60574 0 FreeSans 320 90 0 0 bandgap_trim[1]
port 34 nsew
flabel metal2 416050 60274 416086 60574 0 FreeSans 320 90 0 0 bandgap_trim[0]
port 35 nsew
flabel metal2 405907 66306 406050 66606 0 FreeSans 320 90 0 0 vbgtc
port 36 nsew
flabel metal2 406227 66246 406370 66546 0 FreeSans 320 90 0 0 vbgsc
port 37 nsew
flabel metal3 464466 21962 464808 22139 0 FreeSans 1600 0 0 0 gpio1_1
port 38 nsew
flabel metal1 458471 28689 458531 28958 0 FreeSans 320 90 0 0 vbg_test_to_gpio1_1[1]
port 39 nsew
flabel metal1 458760 28670 458820 28939 0 FreeSans 320 90 0 0 vbg_test_to_gpio1_1[0]
port 40 nsew
<< end >>
