magic
tech sky130A
magscale 1 2
timestamp 1726771202
<< metal1 >>
rect -10325 7780 -10289 13021
rect -5693 7783 -5657 12971
rect -1061 7793 -1025 12995
rect 1038 8677 1095 9530
rect 1038 8620 3095 8677
rect 4725 8641 4761 13997
rect 3038 7653 3095 8620
rect 3571 8605 4761 8641
rect 6015 8690 6072 9561
rect 6015 8633 7727 8690
rect 9721 8649 9757 13889
rect 3571 7783 3607 8605
rect 7670 7614 7727 8633
rect 8203 8613 9757 8649
rect 10992 8658 11049 9528
rect 8203 7792 8239 8613
rect 10992 8601 12359 8658
rect 14667 8631 14703 13857
rect 12302 7641 12359 8601
rect 12835 8595 14703 8631
rect 15969 8654 16026 9570
rect 19629 8663 19665 13915
rect 16934 8654 16991 8659
rect 15969 8597 16991 8654
rect 12835 7788 12871 8595
rect 16934 7648 16991 8597
rect 17467 8627 19665 8663
rect 20946 8662 21003 9545
rect 24533 8677 24569 13953
rect 17467 7779 17503 8627
rect 20946 8605 21623 8662
rect 21566 7643 21623 8605
rect 22099 8641 24569 8677
rect 24653 8684 24689 13957
rect 25639 8684 25645 8697
rect 24653 8648 25645 8684
rect 25639 8645 25645 8648
rect 25697 8645 25703 8697
rect 22099 7993 22135 8641
rect 25923 8192 25980 9615
rect 26723 8645 26729 8697
rect 26781 8645 26787 8697
rect 25923 8135 26257 8192
rect 26198 7644 26255 8135
rect 26735 7987 26771 8645
rect -10858 4375 -10801 5551
rect -6226 4375 -6169 5551
rect -1594 4375 -1537 5551
rect 3038 4375 3095 5551
rect 7670 4375 7727 5551
rect 12302 4375 12359 5551
rect 16934 4375 16991 5551
rect 21566 4375 21623 5551
rect 26198 4375 26255 5545
rect -10863 4367 -10715 4375
rect -10863 4209 -10853 4367
rect -10725 4209 -10715 4367
rect -10863 4197 -10715 4209
rect -6231 4367 -6083 4375
rect -6231 4209 -6221 4367
rect -6093 4209 -6083 4367
rect -6231 4197 -6083 4209
rect -1599 4367 -1451 4375
rect -1599 4209 -1589 4367
rect -1461 4209 -1451 4367
rect -1599 4197 -1451 4209
rect 3033 4367 3181 4375
rect 3033 4209 3043 4367
rect 3171 4209 3181 4367
rect 3033 4197 3181 4209
rect 7665 4367 7813 4375
rect 7665 4209 7675 4367
rect 7803 4209 7813 4367
rect 7665 4197 7813 4209
rect 12297 4367 12445 4375
rect 12297 4209 12307 4367
rect 12435 4209 12445 4367
rect 12297 4197 12445 4209
rect 16929 4367 17077 4375
rect 16929 4209 16939 4367
rect 17067 4209 17077 4367
rect 16929 4197 17077 4209
rect 21561 4367 21709 4375
rect 21561 4209 21571 4367
rect 21699 4209 21709 4367
rect 21561 4197 21709 4209
rect 26193 4367 26341 4375
rect 26193 4209 26203 4367
rect 26331 4209 26341 4367
rect 26193 4197 26341 4209
<< via1 >>
rect 25645 8645 25697 8697
rect 26729 8645 26781 8697
rect -10853 4209 -10725 4367
rect -6221 4209 -6093 4367
rect -1589 4209 -1461 4367
rect 3043 4209 3171 4367
rect 7675 4209 7803 4367
rect 12307 4209 12435 4367
rect 16939 4209 17067 4367
rect 21571 4209 21699 4367
rect 26203 4209 26331 4367
<< metal2 >>
rect 1789 9389 2193 9489
rect 1789 9353 2199 9389
rect -8625 8988 -8196 8991
rect -9192 7591 -8760 8735
rect -8628 7602 -8196 8988
rect -8628 7591 -8620 7602
rect -8204 7591 -8196 7602
rect -4560 7588 -4128 8223
rect -3996 7609 -3564 8465
rect 72 7595 504 7721
rect 636 7608 1068 7975
rect 2027 7018 2199 9353
rect 2378 8541 2573 9353
rect 4045 8892 4240 9371
rect 5848 8892 6016 8893
rect 4045 8697 6016 8892
rect 2378 8352 4556 8541
rect 2398 8351 4556 8352
rect 4366 7989 4556 8351
rect 5848 7989 6016 8697
rect 6655 7018 6827 9401
rect 7355 8541 7550 9421
rect 9022 8924 9217 9403
rect 10480 8924 10648 8925
rect 9022 8729 10648 8924
rect 7352 8351 9188 8541
rect 8998 7989 9188 8351
rect 10480 7989 10648 8729
rect 11291 7018 11463 9397
rect 12332 8541 12527 9381
rect 13999 8908 14194 9387
rect 13999 8903 15218 8908
rect 13999 8713 15280 8903
rect 12332 8354 13820 8541
rect 12348 8351 13820 8354
rect 13630 7989 13820 8351
rect 15112 7989 15280 8713
rect -11788 7015 -11695 7018
rect -7156 7015 -7063 7018
rect -2524 7015 -2431 7018
rect -11869 4425 -11695 7015
rect -11869 3357 -11693 4425
rect -10863 4367 -10715 4375
rect -10863 4209 -10853 4367
rect -10725 4209 -10715 4367
rect -10863 3059 -10715 4209
rect -9530 3639 -9340 4679
rect -8048 3937 -7880 4828
rect -7237 4425 -7063 7015
rect -7237 3357 -7061 4425
rect -6231 4367 -6083 4375
rect -6231 4209 -6221 4367
rect -6093 4209 -6083 4367
rect -6231 3059 -6083 4209
rect -4898 3639 -4708 4679
rect -3416 3937 -3248 4828
rect -2605 4425 -2431 7015
rect -2605 3357 -2429 4425
rect -1599 4367 -1451 4375
rect -1599 4209 -1589 4367
rect -1461 4209 -1451 4367
rect -1599 3059 -1451 4209
rect -266 3639 -76 4679
rect 1216 3937 1384 4828
rect 2027 4425 2201 7018
rect 6655 7003 6833 7018
rect 2027 3357 2203 4425
rect 3033 4367 3181 4375
rect 3033 4209 3043 4367
rect 3171 4209 3181 4367
rect 3033 3059 3181 4209
rect 4366 3639 4556 4679
rect 5848 3937 6016 4828
rect 6659 4425 6833 7003
rect 6659 3357 6835 4425
rect 7665 4367 7813 4375
rect 7665 4209 7675 4367
rect 7803 4209 7813 4367
rect 7665 3059 7813 4209
rect 8998 3639 9188 4679
rect 10480 3937 10648 4828
rect 11291 4425 11465 7018
rect 15925 7015 16097 9383
rect 17309 8617 17504 9375
rect 18976 8641 19171 9403
rect 17309 8422 18452 8617
rect 18976 8541 19908 8641
rect 18976 8446 19912 8541
rect 18262 7989 18452 8422
rect 19744 7989 19912 8446
rect 11291 3357 11467 4425
rect 12297 4367 12445 4375
rect 12297 4209 12307 4367
rect 12435 4209 12445 4367
rect 12297 3059 12445 4209
rect 13630 3639 13820 4679
rect 15112 3937 15280 4828
rect 15923 4425 16097 7015
rect 20553 7018 20725 9375
rect 22286 8587 22481 9363
rect 22286 8392 23084 8587
rect 22894 7989 23084 8392
rect 23953 8555 24148 9391
rect 23953 8360 24544 8555
rect 24376 7989 24544 8360
rect 20553 6977 20729 7018
rect 15923 3357 16099 4425
rect 16929 4367 17077 4375
rect 16929 4209 16939 4367
rect 17067 4209 17077 4367
rect 16929 3059 17077 4209
rect 18262 3639 18452 4679
rect 19744 3937 19912 4828
rect 20555 4425 20729 6977
rect 20555 3357 20731 4425
rect 21561 4367 21709 4375
rect 21561 4209 21571 4367
rect 21699 4209 21709 4367
rect 21561 3059 21709 4209
rect 22894 3639 23084 4679
rect 24376 3937 24544 4828
rect 25187 3357 25363 9374
rect 25645 8697 25697 8703
rect 26729 8697 26781 8703
rect 25697 8653 26729 8689
rect 25645 8639 25697 8645
rect 26729 8639 26781 8645
rect 27263 8615 27458 9391
rect 27263 8420 27716 8615
rect 27526 7989 27716 8420
rect 28930 8541 29125 9379
rect 28930 8310 29176 8541
rect 29008 7989 29176 8310
rect 26193 4367 26341 4375
rect 26193 4209 26203 4367
rect 26331 4209 26341 4367
rect 26193 3059 26341 4209
rect 27526 3639 27716 4529
rect 29008 3937 29176 4551
<< metal3 >>
rect 3697 12950 29596 13080
rect -12973 12694 2902 12824
rect 8685 12438 29596 12568
rect -12973 12182 7890 12312
rect 13660 11926 29596 12056
rect -12973 11670 12851 11800
rect 18652 11414 29596 11544
rect -12973 11158 17848 11288
rect 23563 10902 29596 11032
rect -12973 10646 22832 10776
rect 28578 10390 29596 10520
rect -12973 10134 27829 10264
rect -8580 8854 29596 8984
rect -12973 8598 -8783 8728
rect -3994 8342 29596 8472
rect -12973 8086 -4155 8216
rect 683 7830 29596 7960
rect -12973 7574 477 7704
rect 5364 7318 29596 7448
rect -12973 7062 5058 7192
rect 9959 6806 29596 6936
rect -12973 6550 9708 6680
rect 14572 6294 29596 6424
rect -12973 6038 14340 6168
rect 19217 5782 29596 5912
rect -12973 5526 18990 5656
rect 23840 5270 29596 5400
rect -12973 5014 23609 5144
rect 28482 4758 29596 4888
rect -12973 4502 28236 4632
rect -11993 3955 29595 4155
rect -11993 3655 29595 3855
rect -11993 3355 29595 3555
rect -11993 3055 29595 3255
use cv3_via2_3cut  cv3_via2_3cut_0
timestamp 1719174692
transform 1 0 -538470 0 1 -60112
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_1
timestamp 1719174692
transform 1 0 -532205 0 1 -66261
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_2
timestamp 1719174692
transform 1 0 -513575 0 1 -62670
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_3
timestamp 1719174692
transform 1 0 -519665 0 1 -62425
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_4
timestamp 1719174692
transform 1 0 -518558 0 1 -62154
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_5
timestamp 1719174692
transform 1 0 -524649 0 1 -61898
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_6
timestamp 1719174692
transform 1 0 -523523 0 1 -61637
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_7
timestamp 1719174692
transform 1 0 -529638 0 1 -61395
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_8
timestamp 1719174692
transform 1 0 -528516 0 1 -61139
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_9
timestamp 1719174692
transform 1 0 -534612 0 1 -60873
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_10
timestamp 1719174692
transform 1 0 -533486 0 1 -60622
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_11
timestamp 1719174692
transform 1 0 -539591 0 1 -60366
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_12
timestamp 1719174692
transform 1 0 -514694 0 1 -62926
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_13
timestamp 1719174692
transform 1 0 -514261 0 1 -68554
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_14
timestamp 1719174692
transform 1 0 -513704 0 1 -68307
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_15
timestamp 1719174692
transform 1 0 -518897 0 1 -68050
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_16
timestamp 1719174692
transform 1 0 -518329 0 1 -67793
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_17
timestamp 1719174692
transform 1 0 -523512 0 1 -67536
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_18
timestamp 1719174692
transform 1 0 -522950 0 1 -67279
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_19
timestamp 1719174692
transform 1 0 -528167 0 1 -67022
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_20
timestamp 1719174692
transform 1 0 -527595 0 1 -66760
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_21
timestamp 1719174692
transform 1 0 -532797 0 1 -66494
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_22
timestamp 1719174692
transform 1 0 -550751 0 1 -64210
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_23
timestamp 1719174692
transform 1 0 -537437 0 1 -65990
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_24
timestamp 1719174692
transform 1 0 -536807 0 1 -65742
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_25
timestamp 1719174692
transform 1 0 -542043 0 1 -65476
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_26
timestamp 1719174692
transform 1 0 -541490 0 1 -65219
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_27
timestamp 1719174692
transform 1 0 -546649 0 1 -64967
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_28
timestamp 1719174692
transform 1 0 -546130 0 1 -64729
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_29
timestamp 1719174692
transform 1 0 -551289 0 1 -64467
box 542198 73062 542469 73190
use cv3_via2_8cut  cv3_via2_8cut_0
timestamp 1719106786
transform 0 -1 50671 1 0 -3471
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_1
timestamp 1719106786
transform 0 -1 54331 1 0 -2879
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_2
timestamp 1719106786
transform 0 -1 53013 1 0 -3171
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_3
timestamp 1719106786
transform 0 -1 51485 1 0 -3797
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_4
timestamp 1719106786
transform 0 -1 87727 1 0 -3471
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_5
timestamp 1719106786
transform 0 -1 88541 1 0 -3797
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_6
timestamp 1719106786
transform 0 -1 90069 1 0 -3171
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_7
timestamp 1719106786
transform 0 -1 91387 1 0 -2879
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_8
timestamp 1719106786
transform 0 -1 86755 1 0 -2879
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_9
timestamp 1719106786
transform 0 -1 85437 1 0 -3171
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_10
timestamp 1719106786
transform 0 -1 83909 1 0 -3797
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_11
timestamp 1719106786
transform 0 -1 83095 1 0 -3471
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_12
timestamp 1719106786
transform 0 -1 78463 1 0 -3471
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_13
timestamp 1719106786
transform 0 -1 79277 1 0 -3797
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_14
timestamp 1719106786
transform 0 -1 82123 1 0 -2879
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_15
timestamp 1719106786
transform 0 -1 80805 1 0 -3171
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_16
timestamp 1719106786
transform 0 -1 74645 1 0 -3797
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_17
timestamp 1719106786
transform 0 -1 73831 1 0 -3471
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_18
timestamp 1719106786
transform 0 -1 76173 1 0 -3171
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_19
timestamp 1719106786
transform 0 -1 77491 1 0 -2879
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_20
timestamp 1719106786
transform 0 -1 70013 1 0 -3797
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_21
timestamp 1719106786
transform 0 -1 69199 1 0 -3471
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_22
timestamp 1719106786
transform 0 -1 72859 1 0 -2879
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_23
timestamp 1719106786
transform 0 -1 71541 1 0 -3171
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_24
timestamp 1719106786
transform 0 -1 68227 1 0 -2879
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_25
timestamp 1719106786
transform 0 -1 66909 1 0 -3171
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_26
timestamp 1719106786
transform 0 -1 65381 1 0 -3797
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_27
timestamp 1719106786
transform 0 -1 64567 1 0 -3471
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_28
timestamp 1719106786
transform 0 -1 62277 1 0 -3171
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_29
timestamp 1719106786
transform 0 -1 60749 1 0 -3797
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_30
timestamp 1719106786
transform 0 -1 59935 1 0 -3471
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_31
timestamp 1719106786
transform 0 -1 63595 1 0 -2879
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_32
timestamp 1719106786
transform 0 -1 57645 1 0 -3171
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_33
timestamp 1719106786
transform 0 -1 56117 1 0 -3797
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_34
timestamp 1719106786
transform 0 -1 55303 1 0 -3471
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_35
timestamp 1719106786
transform 0 -1 58963 1 0 -2879
box 6850 62208 6998 62544
use isolated_switch_large  isolated_switch_large_0 ../ip/sky130_ef_ip__analog_switches/mag
array 0 0 4826 0 5 -4977
timestamp 1724442075
transform 0 -1 1366 -1 0 14607
box 660 -3110 5544 1338
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_1 ../ip/sky130_ef_ip__analog_switches/mag
array 0 0 -3542 0 8 -4632
timestamp 1724439637
transform 0 -1 -8220 -1 0 8019
box -4 -600 3538 3648
<< labels >>
flabel metal3 s -12386 4565 -12386 4565 0 FreeSans 960 0 0 0 voutref
flabel metal3 s -12370 5081 -12370 5081 0 FreeSans 960 0 0 0 vinref
flabel metal3 s -12362 5585 -12362 5585 0 FreeSans 960 0 0 0 left_vref
flabel metal3 s -12370 6091 -12370 6091 0 FreeSans 960 0 0 0 right_vref
flabel metal3 s -12434 8155 -12434 8155 0 FreeSans 960 0 0 0 vbgtc
flabel metal3 s -12440 8661 -12440 8661 0 FreeSans 960 0 0 0 vbgsc
flabel metal3 s -12474 11225 -12474 11225 0 FreeSans 960 0 0 0 comp_n
flabel metal3 s -12498 11757 -12498 11757 0 FreeSans 960 0 0 0 comp_p
flabel metal3 s 29198 4822 29198 4822 0 FreeSans 960 0 0 0 user_voutref
flabel metal3 s 29202 5340 29202 5340 0 FreeSans 960 0 0 0 user_vinref
flabel metal3 s 29194 6352 29194 6352 0 FreeSans 960 0 0 0 user_right_vinref
flabel metal3 s 29194 5842 29194 5842 0 FreeSans 960 0 0 0 user_left_vinref
flabel metal3 s 29196 6870 29196 6870 0 FreeSans 960 0 0 0 user_tempsense
flabel metal3 s 29190 7380 29190 7380 0 FreeSans 960 0 0 0 user_dac0
flabel metal3 s 29198 7904 29198 7904 0 FreeSans 960 0 0 0 user_dac1
flabel metal3 s 29202 8406 29202 8406 0 FreeSans 960 0 0 0 user_vbgtc
flabel metal3 s 29166 8912 29166 8912 0 FreeSans 960 0 0 0 user_vbgsc
flabel metal3 s 29134 10444 29134 10444 0 FreeSans 960 0 0 0 user_adc0
flabel metal3 s 29134 10962 29134 10962 0 FreeSans 960 0 0 0 user_adc1
flabel metal3 s 29132 11480 29132 11480 0 FreeSans 960 0 0 0 user_comp_n
flabel metal3 s 29138 11988 29138 11988 0 FreeSans 960 0 0 0 user_comp_p
flabel metal3 s 29132 12504 29132 12504 0 FreeSans 960 0 0 0 user_ulpcomp_n
flabel metal3 s 29138 13008 29138 13008 0 FreeSans 960 0 0 0 user_ulpcomp_p
flabel metal3 s -12518 12741 -12518 12741 0 FreeSans 960 0 0 0 ulpcomp_p
flabel metal3 s -12508 12249 -12508 12249 0 FreeSans 960 0 0 0 ulpcomp_n
flabel metal3 s -12456 10705 -12456 10705 0 FreeSans 960 0 0 0 adc1
flabel metal3 s -12444 10193 -12444 10193 0 FreeSans 960 0 0 0 adc0
flabel metal3 s -12430 7641 -12430 7641 0 FreeSans 960 0 0 0 dac1
flabel metal3 s -12424 7101 -12424 7101 0 FreeSans 960 0 0 0 dac0
flabel metal3 s -12434 6611 -12434 6611 0 FreeSans 960 0 0 0 tempsense
flabel metal3 s -11306 4056 -11306 4056 0 FreeSans 960 0 0 0 vssa0
flabel metal3 s -11316 3756 -11316 3756 0 FreeSans 960 0 0 0 vdda0
flabel metal3 s -11326 3146 -11326 3146 0 FreeSans 960 0 0 0 vccd0
flabel metal3 s -11306 3462 -11306 3462 0 FreeSans 960 0 0 0 vssd0
<< end >>
