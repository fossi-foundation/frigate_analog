VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_routes_left
  CLASS COVER ;
  FOREIGN analog_routes_left ;
  ORIGIN 0.000 0.000 ;
  SIZE 190.595 BY 2509.385 ;
  OBS
      LAYER met2 ;
        RECT -1.280 1468.955 -1.040 1480.495 ;
        RECT -1.280 1304.115 -1.040 1315.345 ;
        RECT -1.280 1139.045 -1.040 1150.295 ;
        RECT -1.280 961.115 -1.040 985.385 ;
        RECT -1.280 960.875 -0.145 961.115 ;
        RECT -0.385 851.065 -0.145 960.875 ;
        RECT 0.975 851.065 2.245 851.725 ;
        RECT -1.865 850.825 2.245 851.065 ;
        RECT 0.975 850.475 2.245 850.825 ;
        RECT -0.585 800.215 0.795 800.455 ;
        RECT 0.555 660.715 0.795 800.215 ;
        RECT -1.280 660.475 0.795 660.715 ;
        RECT -1.280 651.135 -1.040 660.475 ;
        RECT -1.280 486.135 -1.040 497.175 ;
        RECT -1.280 321.055 -1.040 332.145 ;
        RECT -1.280 156.055 -1.040 167.315 ;
      LAYER met3 ;
        RECT 1.210 2450.985 4.710 2451.625 ;
        RECT 1.210 2345.985 4.710 2346.625 ;
        RECT 1.210 2240.985 4.710 2241.625 ;
        RECT 1.210 2135.985 4.710 2136.625 ;
        RECT 1.210 1482.735 4.710 1482.775 ;
        RECT 0.000 1482.135 4.710 1482.735 ;
        RECT 1.210 1317.735 4.710 1317.775 ;
        RECT 0.000 1317.135 4.710 1317.735 ;
        RECT 1.210 1152.735 4.710 1152.775 ;
        RECT 0.000 1152.135 4.710 1152.735 ;
        RECT 1.210 987.735 4.710 987.775 ;
        RECT 0.000 987.135 4.710 987.735 ;
        RECT 2.855 852.010 4.355 852.155 ;
        RECT 1.315 851.725 4.355 852.010 ;
        RECT 0.975 850.475 4.355 851.725 ;
        RECT 1.315 850.010 4.355 850.475 ;
        RECT 2.855 848.025 4.355 850.010 ;
        RECT 1.210 800.020 4.710 800.660 ;
        RECT 1.210 499.735 4.710 499.775 ;
        RECT 1.205 499.135 4.710 499.735 ;
        RECT 1.210 334.735 4.710 334.775 ;
        RECT 0.000 334.135 4.710 334.735 ;
        RECT 1.210 171.020 4.710 171.060 ;
        RECT 0.000 170.420 4.710 171.020 ;
        RECT 1.210 6.020 4.710 6.060 ;
        RECT 0.000 5.420 4.710 6.020 ;
      LAYER met4 ;
        RECT 156.635 2457.165 157.275 2509.385 ;
        RECT 154.070 2455.565 157.275 2457.165 ;
        RECT 156.635 2455.560 157.275 2455.565 ;
        RECT 157.935 2452.165 158.575 2509.385 ;
        RECT 2.260 2451.625 4.740 2452.165 ;
        RECT 1.210 2450.985 4.740 2451.625 ;
        RECT 2.260 2450.565 4.740 2450.985 ;
        RECT 155.375 2450.565 158.575 2452.165 ;
        RECT 159.195 2447.165 159.835 2509.385 ;
        RECT 156.635 2445.565 159.835 2447.165 ;
        RECT 159.195 2352.165 159.835 2445.565 ;
        RECT 156.630 2350.565 159.835 2352.165 ;
        RECT 159.195 2350.555 159.835 2350.565 ;
        RECT 160.495 2347.165 161.135 2509.385 ;
        RECT 2.260 2346.625 4.740 2347.165 ;
        RECT 1.210 2345.985 4.740 2346.625 ;
        RECT 2.260 2345.565 4.740 2345.985 ;
        RECT 157.940 2345.565 161.140 2347.165 ;
        RECT 161.755 2342.165 162.395 2509.385 ;
        RECT 159.195 2340.565 162.395 2342.165 ;
        RECT 161.755 2247.170 162.395 2340.565 ;
        RECT 159.195 2245.570 162.395 2247.170 ;
        RECT 161.755 2245.560 162.395 2245.570 ;
        RECT 163.055 2242.165 163.695 2509.385 ;
        RECT 2.260 2241.625 4.740 2242.165 ;
        RECT 1.210 2240.985 4.740 2241.625 ;
        RECT 2.260 2240.565 4.740 2240.985 ;
        RECT 160.495 2240.565 163.695 2242.165 ;
        RECT 164.315 2237.160 164.955 2509.385 ;
        RECT 161.750 2235.560 164.955 2237.160 ;
        RECT 164.315 2142.165 164.955 2235.560 ;
        RECT 161.755 2140.565 164.955 2142.165 ;
        RECT 164.315 2140.515 164.955 2140.565 ;
        RECT 165.615 2137.165 166.255 2509.385 ;
        RECT 2.260 2136.625 4.740 2137.165 ;
        RECT 1.210 2135.985 4.740 2136.625 ;
        RECT 2.260 2135.565 4.740 2135.985 ;
        RECT 163.060 2135.565 166.260 2137.165 ;
        RECT 166.875 2132.175 167.515 2509.385 ;
        RECT 164.320 2130.575 167.520 2132.175 ;
        RECT 166.875 1488.305 167.515 2130.575 ;
        RECT 164.315 1486.705 167.515 1488.305 ;
        RECT 168.175 1483.325 168.815 2509.385 ;
        RECT 2.260 1482.775 4.740 1483.320 ;
        RECT 1.210 1482.135 4.740 1482.775 ;
        RECT 2.260 1481.715 4.740 1482.135 ;
        RECT 165.615 1481.725 168.815 1483.325 ;
        RECT 169.435 1478.305 170.075 2509.385 ;
        RECT 166.880 1476.705 170.080 1478.305 ;
        RECT 169.435 1323.300 170.075 1476.705 ;
        RECT 166.880 1321.700 170.080 1323.300 ;
        RECT 169.435 1321.680 170.075 1321.700 ;
        RECT 2.260 1317.775 4.740 1318.315 ;
        RECT 170.735 1318.295 171.375 2509.385 ;
        RECT 1.210 1317.135 4.740 1317.775 ;
        RECT 2.260 1316.715 4.740 1317.135 ;
        RECT 168.175 1316.695 171.375 1318.295 ;
        RECT 171.995 1313.305 172.635 2509.385 ;
        RECT 169.435 1311.705 172.635 1313.305 ;
        RECT 171.995 1158.425 172.635 1311.705 ;
        RECT 169.440 1156.825 172.640 1158.425 ;
        RECT 171.995 1156.805 172.635 1156.825 ;
        RECT 173.295 1153.435 173.935 2509.385 ;
        RECT 2.260 1152.775 4.740 1153.315 ;
        RECT 1.210 1152.135 4.740 1152.775 ;
        RECT 2.260 1151.715 4.740 1152.135 ;
        RECT 170.735 1151.835 173.935 1153.435 ;
        RECT 174.555 1148.440 175.195 2509.385 ;
        RECT 172.000 1146.840 175.200 1148.440 ;
        RECT 174.555 993.300 175.195 1146.840 ;
        RECT 171.995 991.700 175.195 993.300 ;
        RECT 2.260 987.775 4.740 988.315 ;
        RECT 175.855 988.310 176.495 2509.385 ;
        RECT 1.210 987.135 4.740 987.775 ;
        RECT 2.260 986.715 4.740 987.135 ;
        RECT 173.295 986.710 176.495 988.310 ;
        RECT 177.115 983.305 177.755 2509.385 ;
        RECT 174.565 981.705 177.765 983.305 ;
        RECT 2.855 848.025 4.355 852.155 ;
        RECT 3.225 801.200 3.985 848.025 ;
        RECT 177.115 806.205 177.755 981.705 ;
        RECT 174.555 804.605 177.755 806.205 ;
        RECT 177.115 804.595 177.755 804.605 ;
        RECT 178.415 801.200 179.055 2509.385 ;
        RECT 2.260 800.660 4.740 801.200 ;
        RECT 1.210 800.020 4.740 800.660 ;
        RECT 2.260 799.600 4.740 800.020 ;
        RECT 175.855 799.600 179.055 801.200 ;
        RECT 179.675 796.205 180.315 2509.385 ;
        RECT 177.110 794.605 180.315 796.205 ;
        RECT 179.675 505.300 180.315 794.605 ;
        RECT 177.115 503.700 180.315 505.300 ;
        RECT 2.260 499.775 4.740 500.315 ;
        RECT 180.975 500.310 181.615 2509.385 ;
        RECT 1.210 499.135 4.740 499.775 ;
        RECT 2.260 498.715 4.740 499.135 ;
        RECT 178.425 498.710 181.625 500.310 ;
        RECT 182.235 495.310 182.875 2509.385 ;
        RECT 179.675 493.710 182.875 495.310 ;
        RECT 182.235 340.295 182.875 493.710 ;
        RECT 179.665 338.705 182.875 340.295 ;
        RECT 179.665 338.695 182.865 338.705 ;
        RECT 2.260 334.775 4.740 335.315 ;
        RECT 183.535 335.295 184.175 2509.385 ;
        RECT 1.210 334.135 4.740 334.775 ;
        RECT 2.260 333.715 4.740 334.135 ;
        RECT 180.975 333.695 184.175 335.295 ;
        RECT 184.795 330.295 185.435 2509.385 ;
        RECT 182.235 328.695 185.435 330.295 ;
        RECT 184.795 176.605 185.435 328.695 ;
        RECT 182.235 175.005 185.435 176.605 ;
        RECT 2.260 171.060 4.740 171.600 ;
        RECT 186.095 171.575 186.735 2509.385 ;
        RECT 1.210 170.420 4.740 171.060 ;
        RECT 2.260 170.000 4.740 170.420 ;
        RECT 183.535 169.975 186.735 171.575 ;
        RECT 187.355 166.605 187.995 2509.385 ;
        RECT 184.800 165.005 188.000 166.605 ;
        RECT 187.355 11.575 187.995 165.005 ;
        RECT 184.675 9.975 187.995 11.575 ;
        RECT 187.355 9.935 187.995 9.975 ;
        RECT 2.260 6.060 4.740 6.600 ;
        RECT 188.655 6.595 189.295 2509.385 ;
        RECT 1.210 5.420 4.740 6.060 ;
        RECT 2.260 5.000 4.740 5.420 ;
        RECT 186.095 4.995 189.295 6.595 ;
        RECT 189.955 1.720 190.595 2509.385 ;
        RECT 187.275 0.120 190.595 1.720 ;
        RECT 189.955 0.000 190.595 0.120 ;
      LAYER met5 ;
        RECT 153.950 2457.165 157.390 2457.285 ;
        RECT 4.620 2455.565 157.455 2457.165 ;
        RECT 153.950 2455.445 157.390 2455.565 ;
        RECT 155.255 2452.165 158.695 2452.285 ;
        RECT 2.260 2450.565 158.695 2452.165 ;
        RECT 155.255 2450.445 158.695 2450.565 ;
        RECT 156.515 2447.165 159.955 2447.285 ;
        RECT 4.620 2445.565 159.955 2447.165 ;
        RECT 156.515 2445.445 159.955 2445.565 ;
        RECT 156.510 2352.165 159.950 2352.285 ;
        RECT 4.620 2350.565 160.015 2352.165 ;
        RECT 156.510 2350.445 159.950 2350.565 ;
        RECT 157.820 2347.165 161.260 2347.285 ;
        RECT 2.260 2345.565 161.260 2347.165 ;
        RECT 157.820 2345.445 161.260 2345.565 ;
        RECT 159.075 2342.165 162.515 2342.285 ;
        RECT 4.620 2340.565 162.515 2342.165 ;
        RECT 159.075 2340.445 162.515 2340.565 ;
        RECT 159.075 2247.165 162.515 2247.290 ;
        RECT 4.620 2245.565 162.575 2247.165 ;
        RECT 159.075 2245.450 162.515 2245.565 ;
        RECT 160.375 2242.165 163.815 2242.285 ;
        RECT 2.260 2240.565 163.815 2242.165 ;
        RECT 160.375 2240.445 163.815 2240.565 ;
        RECT 161.630 2237.165 165.070 2237.280 ;
        RECT 4.620 2235.565 165.070 2237.165 ;
        RECT 161.630 2235.440 165.070 2235.565 ;
        RECT 161.635 2142.165 165.075 2142.285 ;
        RECT 4.620 2140.565 165.135 2142.165 ;
        RECT 161.635 2140.445 165.075 2140.565 ;
        RECT 162.940 2137.165 166.380 2137.285 ;
        RECT 2.260 2135.565 166.380 2137.165 ;
        RECT 162.940 2135.445 166.380 2135.565 ;
        RECT 164.200 2132.165 167.640 2132.295 ;
        RECT 4.620 2130.565 167.640 2132.165 ;
        RECT 164.200 2130.455 167.640 2130.565 ;
        RECT 164.195 1488.320 167.635 1488.425 ;
        RECT 4.620 1486.720 167.695 1488.320 ;
        RECT 164.195 1486.585 167.635 1486.720 ;
        RECT 165.495 1483.320 168.935 1483.445 ;
        RECT 2.260 1481.720 168.935 1483.320 ;
        RECT 165.495 1481.605 168.935 1481.720 ;
        RECT 166.760 1478.320 170.200 1478.425 ;
        RECT 4.620 1476.720 170.200 1478.320 ;
        RECT 166.760 1476.585 170.200 1476.720 ;
        RECT 166.760 1323.315 170.200 1323.420 ;
        RECT 4.620 1321.715 170.255 1323.315 ;
        RECT 166.760 1321.580 170.200 1321.715 ;
        RECT 168.055 1318.315 171.495 1318.415 ;
        RECT 2.260 1316.715 171.495 1318.315 ;
        RECT 168.055 1316.575 171.495 1316.715 ;
        RECT 169.315 1313.315 172.755 1313.425 ;
        RECT 4.620 1311.715 172.755 1313.315 ;
        RECT 169.315 1311.585 172.755 1311.715 ;
        RECT 169.320 1158.450 172.760 1158.545 ;
        RECT 4.620 1156.850 172.815 1158.450 ;
        RECT 169.320 1156.705 172.760 1156.850 ;
        RECT 170.615 1153.450 174.055 1153.555 ;
        RECT 3.015 1153.315 174.055 1153.450 ;
        RECT 2.260 1151.850 174.055 1153.315 ;
        RECT 2.260 1151.715 5.065 1151.850 ;
        RECT 170.615 1151.715 174.055 1151.850 ;
        RECT 171.880 1148.450 175.320 1148.560 ;
        RECT 4.620 1146.850 175.320 1148.450 ;
        RECT 171.880 1146.720 175.320 1146.850 ;
        RECT 171.875 993.315 175.315 993.420 ;
        RECT 4.620 991.715 175.375 993.315 ;
        RECT 171.875 991.580 175.315 991.715 ;
        RECT 173.175 988.315 176.615 988.430 ;
        RECT 2.260 986.715 176.615 988.315 ;
        RECT 173.175 986.590 176.615 986.715 ;
        RECT 174.445 983.315 177.885 983.425 ;
        RECT 4.620 981.715 177.885 983.315 ;
        RECT 174.445 981.585 177.885 981.715 ;
        RECT 174.435 806.200 177.875 806.325 ;
        RECT 4.620 804.600 177.935 806.200 ;
        RECT 174.435 804.485 177.875 804.600 ;
        RECT 175.735 801.200 179.175 801.320 ;
        RECT 2.260 799.600 179.175 801.200 ;
        RECT 175.735 799.480 179.175 799.600 ;
        RECT 176.990 796.200 180.430 796.325 ;
        RECT 4.620 794.600 180.430 796.200 ;
        RECT 176.990 794.485 180.430 794.600 ;
        RECT 176.995 505.315 180.435 505.420 ;
        RECT 4.620 503.715 180.495 505.315 ;
        RECT 176.995 503.580 180.435 503.715 ;
        RECT 178.305 500.315 181.745 500.430 ;
        RECT 2.260 498.715 181.745 500.315 ;
        RECT 178.305 498.590 181.745 498.715 ;
        RECT 179.555 495.315 182.995 495.430 ;
        RECT 4.620 493.715 182.995 495.315 ;
        RECT 179.555 493.590 182.995 493.715 ;
        RECT 179.545 340.315 182.985 340.415 ;
        RECT 4.620 338.715 183.055 340.315 ;
        RECT 179.545 338.575 182.985 338.715 ;
        RECT 180.855 335.315 184.295 335.415 ;
        RECT 2.260 333.715 184.295 335.315 ;
        RECT 180.855 333.575 184.295 333.715 ;
        RECT 182.115 330.315 185.555 330.415 ;
        RECT 4.620 328.715 185.555 330.315 ;
        RECT 182.115 328.575 185.555 328.715 ;
        RECT 182.115 176.600 185.555 176.725 ;
        RECT 4.620 175.000 185.555 176.600 ;
        RECT 182.115 174.885 185.555 175.000 ;
        RECT 183.415 171.600 186.855 171.695 ;
        RECT 2.260 170.000 186.855 171.600 ;
        RECT 183.415 169.855 186.855 170.000 ;
        RECT 184.680 166.600 188.120 166.725 ;
        RECT 4.620 165.000 188.120 166.600 ;
        RECT 184.680 164.885 188.120 165.000 ;
        RECT 184.555 11.600 187.995 11.695 ;
        RECT 4.620 10.000 188.175 11.600 ;
        RECT 184.555 9.855 187.995 10.000 ;
        RECT 185.975 6.600 189.415 6.715 ;
        RECT 2.260 5.000 189.415 6.600 ;
        RECT 185.975 4.875 189.415 5.000 ;
        RECT 187.155 1.600 190.595 1.840 ;
        RECT 4.620 0.000 190.595 1.600 ;
  END
END analog_routes_left
END LIBRARY

