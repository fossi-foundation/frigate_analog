magic
tech sky130A
magscale 1 2
timestamp 1738189644
<< checkpaint >>
rect 13576 90470 44674 108774
rect 11788 89638 44674 90470
rect 11788 77304 24064 89638
rect 47564 79666 51798 106318
rect 90466 101676 103632 102450
rect 90370 90174 103632 101676
rect 170731 88410 174936 106921
rect 179684 88392 183889 106903
rect 286916 104224 294176 104230
rect 286916 103456 312116 104224
rect 266368 102290 279534 103064
rect 266272 90788 279534 102290
rect 11788 77208 23290 77304
rect 142418 77026 157512 83794
rect 160821 80030 176451 87002
rect 178169 80012 193799 86984
rect 211561 84325 214208 85072
rect 211561 84082 214983 84325
rect 211561 83930 215241 84082
rect 286820 83936 312116 103456
rect 314970 102038 328136 102812
rect 314874 90536 328136 102038
rect 405109 87958 409314 106469
rect 413762 87898 417967 106409
rect 492258 102000 505424 102774
rect 492258 90498 505520 102000
rect 197980 83912 215241 83930
rect 197980 79561 229414 83912
rect 197980 79541 214208 79561
rect 197980 77162 213074 79541
rect 214320 77144 229414 79561
rect 230320 77144 245414 83912
rect 292916 75876 312116 83936
rect 375164 77156 390258 83924
rect 395199 79578 410829 86550
rect 412247 79518 427877 86490
rect 434754 77222 449848 83990
rect 453196 77324 472806 84092
rect 476596 77324 496206 84092
rect 509682 82422 513916 109074
rect 551674 82191 563950 95357
rect 551674 82095 563176 82191
rect 201508 73979 204562 73980
rect 30660 71458 204562 73979
rect 364760 70794 385406 76447
rect 387890 70794 408536 76447
rect 411020 70794 431666 76447
rect 434150 70794 454796 76447
rect 457280 70794 473300 76447
rect 475784 70794 487178 76447
rect 489662 70794 501056 76447
rect 364757 64732 505679 70794
rect 11944 49105 24220 62271
rect 11944 49009 23446 49105
rect 11944 35109 24220 48275
rect 11944 35013 23446 35109
rect 11944 20913 24220 34079
rect 11944 20817 23446 20913
rect 36368 14121 80561 56390
rect 83091 22359 89988 36008
rect 125036 22359 131933 36008
rect 90933 9868 106568 17319
rect 108456 9868 124091 17319
rect 133443 7807 171660 61295
rect 177980 53774 183184 57634
rect 186359 51217 192179 55451
rect 174562 27160 178796 32116
rect 192395 7945 230612 61433
rect 236238 51028 282944 62429
rect 254302 41762 282944 51028
rect 341762 45375 347824 57271
rect 362931 48629 374889 59417
rect 483288 58289 522024 62262
rect 546930 61534 567594 81141
rect 401943 45565 405647 49725
rect 231982 27328 236216 32284
rect 272928 32028 276388 32124
rect 272928 18862 277162 32028
rect 341762 13522 353748 45375
rect 382030 39919 386264 45381
rect 416229 45288 422049 48953
rect 371322 20029 386320 39919
rect 391895 20266 431718 45288
rect 435584 20672 453516 43758
rect 341762 13447 347824 13522
rect 133512 6692 171588 7807
rect 192464 6830 230540 7945
rect 362312 6040 409736 17423
rect 483242 16155 522024 58289
rect 529471 56206 542733 59666
rect 529567 55432 542733 56206
rect 530855 34809 535089 47975
rect 543824 47874 556100 61040
rect 543824 47803 555326 47874
rect 542974 47778 555326 47803
rect 530855 34713 534315 34809
rect 542974 34637 555250 47778
rect 542974 34541 554476 34637
rect 530826 21244 535060 34410
rect 542674 21250 554950 34416
rect 530826 21148 534286 21244
rect 542674 21154 554176 21250
rect 463349 8756 522024 16155
rect 463349 7037 484145 8756
<< error_p >>
rect 77455 38554 77456 38608
rect 77515 38504 77516 38554
rect 77515 38234 77516 38318
<< error_s >>
rect 87646 57219 87648 57881
rect 87700 57219 87702 57881
rect 95783 54285 95785 57546
rect 95837 54241 95839 57502
rect 99327 54610 99329 57895
rect 99381 54610 99383 57895
rect 110361 56992 110365 57026
rect 100583 54502 100617 54525
rect 100583 54464 100655 54487
rect 113479 52688 113490 52756
rect 87646 45301 87648 45963
rect 87700 45301 87702 45963
rect 95783 42367 95785 45628
rect 95837 42323 95839 45584
rect 99327 42692 99329 45977
rect 99381 42692 99383 45977
rect 110361 45074 110365 45108
rect 100583 42584 100617 42607
rect 100583 42546 100655 42569
rect 113479 40819 113490 40838
<< metal1 >>
rect 509660 112322 571519 112362
rect 571571 112322 571586 112362
rect 504650 110336 504656 110388
rect 504708 110382 504714 110388
rect 509660 110382 509700 112322
rect 504708 110342 509700 110382
rect 509780 112202 571399 112242
rect 571451 112202 571468 112242
rect 504708 110336 504714 110342
rect 504530 110216 504536 110268
rect 504588 110262 504594 110268
rect 509780 110262 509820 112202
rect 504588 110222 509820 110262
rect 509900 112082 571279 112122
rect 571331 112082 571344 112122
rect 504588 110216 504594 110222
rect 504890 110096 504896 110148
rect 504948 110142 504954 110148
rect 509900 110142 509940 112082
rect 504948 110102 509940 110142
rect 510020 111962 571159 112002
rect 571211 111962 571218 112002
rect 504948 110096 504954 110102
rect 504768 109976 504774 110028
rect 504826 110022 504832 110028
rect 510020 110022 510060 111962
rect 504826 109982 510060 110022
rect 510140 111842 571039 111882
rect 571091 111842 571098 111882
rect 504826 109976 504832 109982
rect 498982 109902 498988 109908
rect 498968 109862 498988 109902
rect 498982 109856 498988 109862
rect 499040 109902 499046 109908
rect 510140 109902 510180 111842
rect 499040 109862 510180 109902
rect 510260 111722 570919 111762
rect 570971 111722 570990 111762
rect 499040 109856 499046 109862
rect 498870 109782 498876 109788
rect 498850 109742 498876 109782
rect 498870 109736 498876 109742
rect 498928 109782 498934 109788
rect 510260 109782 510300 111722
rect 498928 109742 510300 109782
rect 510380 111602 570799 111642
rect 570851 111602 570870 111642
rect 498928 109736 498934 109742
rect 498740 109662 498746 109668
rect 498710 109622 498746 109662
rect 498740 109616 498746 109622
rect 498798 109662 498804 109668
rect 510380 109662 510420 111602
rect 498798 109622 510420 109662
rect 510500 111482 570679 111522
rect 570731 111482 570748 111522
rect 498798 109616 498804 109622
rect 498620 109542 498626 109548
rect 498604 109502 498626 109542
rect 498620 109496 498626 109502
rect 498678 109542 498684 109548
rect 510500 109542 510540 111482
rect 498678 109502 510540 109542
rect 510620 111362 570559 111402
rect 570611 111362 570624 111402
rect 498678 109496 498684 109502
rect 321590 109376 321596 109428
rect 321648 109422 321654 109428
rect 510620 109422 510660 111362
rect 321648 109382 510660 109422
rect 510740 111242 570439 111282
rect 570491 111242 570506 111282
rect 321648 109376 321654 109382
rect 321712 109256 321718 109308
rect 321770 109302 321776 109308
rect 510740 109302 510780 111242
rect 321770 109262 510780 109302
rect 510860 111122 570319 111162
rect 570371 111122 570386 111162
rect 321770 109256 321776 109262
rect 321344 109136 321350 109188
rect 321402 109182 321408 109188
rect 510860 109182 510900 111122
rect 321402 109142 510900 109182
rect 510980 111002 570199 111042
rect 570251 111002 570266 111042
rect 321402 109136 321408 109142
rect 91299 109059 91305 109069
rect 10603 109027 10606 109059
rect 10658 109027 91305 109059
rect 91299 109017 91305 109027
rect 91357 109059 91363 109069
rect 91357 109027 91377 109059
rect 91357 109017 91363 109027
rect 321462 109016 321468 109068
rect 321520 109062 321526 109068
rect 510980 109062 511020 111002
rect 321520 109022 511020 109062
rect 511100 110882 570079 110922
rect 570131 110882 570140 110922
rect 321520 109016 321526 109022
rect 91176 108987 91182 108997
rect 10760 108955 91182 108987
rect 91176 108945 91182 108955
rect 91234 108987 91240 108997
rect 91234 108955 91252 108987
rect 91234 108945 91240 108955
rect 91046 108915 91052 108925
rect 10873 108883 91052 108915
rect 91046 108873 91052 108883
rect 91104 108873 91110 108925
rect 315440 108896 315446 108948
rect 315498 108942 315504 108948
rect 511100 108942 511140 110882
rect 315498 108902 511140 108942
rect 511220 110762 569959 110802
rect 570011 110762 570024 110802
rect 315498 108896 315504 108902
rect 90930 108843 90936 108853
rect 10941 108840 90936 108843
rect 10987 108811 90936 108840
rect 90930 108801 90936 108811
rect 90988 108801 90994 108853
rect 96959 108771 96965 108781
rect 11045 108766 96965 108771
rect 11097 108739 96965 108766
rect 96959 108729 96965 108739
rect 97017 108771 97023 108781
rect 315552 108776 315558 108828
rect 315610 108822 315616 108828
rect 511220 108822 511260 110762
rect 315610 108782 511260 108822
rect 511340 110642 569841 110682
rect 569893 110642 569902 110682
rect 315610 108776 315616 108782
rect 97017 108739 97036 108771
rect 97017 108729 97023 108739
rect 96840 108699 96846 108709
rect 11204 108667 96846 108699
rect 96840 108657 96846 108667
rect 96898 108699 96904 108709
rect 96898 108667 96921 108699
rect 96898 108657 96904 108667
rect 315672 108656 315678 108708
rect 315730 108702 315736 108708
rect 511340 108702 511380 110642
rect 315730 108662 511380 108702
rect 511460 110522 569717 110562
rect 569769 110522 569790 110562
rect 315730 108656 315736 108662
rect 97202 108627 97208 108637
rect 11322 108595 97208 108627
rect 97202 108585 97208 108595
rect 97260 108627 97266 108637
rect 97260 108595 97273 108627
rect 97260 108585 97266 108595
rect 97078 108555 97084 108565
rect 11424 108523 97084 108555
rect 97078 108513 97084 108523
rect 97136 108555 97142 108565
rect 97136 108523 97148 108555
rect 315798 108536 315804 108588
rect 315856 108582 315862 108588
rect 511460 108582 511500 110522
rect 315856 108542 511500 108582
rect 315856 108536 315862 108542
rect 97136 108513 97142 108523
rect 267209 108489 267261 108495
rect 11718 108477 267209 108479
rect 11766 108447 267209 108477
rect 267261 108447 267270 108479
rect 267209 108431 267261 108437
rect 267083 108407 267089 108417
rect 11874 108375 267089 108407
rect 267083 108365 267089 108375
rect 267141 108407 267147 108417
rect 267141 108375 267149 108407
rect 267141 108365 267147 108375
rect 266958 108335 266964 108345
rect 11941 108330 266964 108335
rect 11990 108303 266964 108330
rect 266958 108293 266964 108303
rect 267016 108335 267022 108345
rect 267016 108303 267027 108335
rect 267016 108293 267022 108303
rect 266834 108263 266840 108273
rect 12096 108231 266840 108263
rect 266834 108221 266840 108231
rect 266892 108263 266898 108273
rect 266892 108231 266900 108263
rect 266892 108221 266898 108231
rect 272866 108191 272872 108201
rect 12218 108159 272872 108191
rect 272866 108149 272872 108159
rect 272924 108191 272930 108201
rect 272924 108159 272936 108191
rect 272924 108149 272930 108159
rect 272741 108119 272747 108129
rect 12277 108087 12280 108119
rect 12332 108087 272747 108119
rect 272741 108077 272747 108087
rect 272799 108119 272805 108129
rect 272799 108087 272818 108119
rect 272799 108077 272805 108087
rect 12385 108042 273155 108047
rect 12385 108015 12389 108042
rect 12441 108015 273155 108042
rect 12503 107968 273034 107975
rect 12551 107943 273034 107968
rect 266834 107819 266840 107871
rect 266892 107819 266898 107871
rect 266850 107744 266882 107819
rect 266957 107816 266963 107868
rect 267015 107816 267021 107868
rect 267085 107854 267137 107860
rect 90936 107729 90988 107735
rect 91053 107686 91059 107738
rect 91111 107686 91117 107738
rect 266973 107735 267005 107816
rect 267204 107812 267210 107864
rect 267262 107812 267268 107864
rect 272741 107840 272747 107892
rect 272799 107840 272805 107892
rect 272866 107849 272872 107901
rect 272924 107849 272930 107901
rect 267085 107737 267137 107802
rect 90936 107671 90988 107677
rect 90946 107115 90978 107671
rect 91069 107122 91101 107686
rect 91176 107670 91182 107722
rect 91234 107670 91240 107722
rect 91292 107677 91298 107729
rect 91350 107677 91356 107729
rect 91192 107117 91224 107670
rect 91308 107115 91340 107677
rect 96840 107659 96846 107711
rect 96898 107659 96904 107711
rect 96856 107126 96888 107659
rect 96959 107647 96965 107699
rect 97017 107647 97023 107699
rect 97078 107668 97084 107720
rect 97136 107668 97142 107720
rect 267220 107716 267252 107812
rect 272757 107704 272789 107840
rect 272882 107739 272914 107849
rect 273002 107737 273034 107943
rect 273123 107744 273155 108015
rect 321718 107950 321770 107956
rect 321344 107886 321350 107938
rect 321402 107886 321408 107938
rect 321462 107886 321468 107938
rect 321520 107886 321526 107938
rect 321590 107896 321596 107948
rect 321648 107896 321654 107948
rect 315440 107710 315446 107762
rect 315498 107710 315504 107762
rect 315550 107720 315556 107772
rect 315608 107720 315614 107772
rect 315672 107734 315678 107786
rect 315730 107734 315736 107786
rect 315798 107734 315804 107786
rect 315856 107734 315862 107786
rect 96975 107135 97007 107647
rect 97094 107135 97126 107668
rect 97202 107647 97208 107699
rect 97260 107647 97266 107699
rect 97218 107123 97250 107647
rect 315452 107458 315492 107710
rect 315562 107448 315602 107720
rect 315684 107450 315724 107734
rect 315810 107432 315850 107734
rect 321356 107448 321396 107886
rect 321474 107472 321514 107886
rect 321602 107478 321642 107896
rect 321718 107892 321770 107898
rect 321724 107454 321764 107892
rect 498620 107818 498626 107870
rect 498678 107818 498684 107870
rect 504536 107860 504588 107866
rect 498632 107436 498672 107818
rect 498740 107806 498746 107858
rect 498798 107806 498804 107858
rect 498870 107808 498876 107860
rect 498928 107808 498934 107860
rect 498752 107416 498792 107806
rect 498882 107410 498922 107808
rect 498982 107806 498988 107858
rect 499040 107806 499046 107858
rect 504650 107818 504656 107870
rect 504708 107818 504714 107870
rect 504768 107830 504774 107882
rect 504826 107830 504832 107882
rect 498994 107414 499034 107806
rect 504536 107802 504588 107808
rect 504542 107420 504582 107802
rect 504662 107420 504702 107818
rect 504780 107416 504820 107830
rect 504890 107828 504896 107880
rect 504948 107828 504954 107880
rect 504902 107430 504942 107828
rect 509044 107360 509080 107370
rect 509025 107354 509105 107360
rect 509025 107268 509105 107274
rect 508950 104952 508986 104961
rect 508926 104946 509006 104952
rect 508926 104860 509006 104866
rect 48461 104556 48497 104566
rect 48440 104550 48520 104556
rect 48440 104464 48520 104470
rect 45394 102586 45400 102594
rect 43378 102550 45400 102586
rect 45394 102542 45400 102550
rect 45452 102586 45458 102594
rect 45452 102550 45463 102586
rect 45452 102542 45458 102550
rect 45310 102502 45316 102510
rect 43378 102466 45316 102502
rect 45310 102458 45316 102466
rect 45368 102502 45374 102510
rect 45368 102466 45384 102502
rect 45368 102458 45374 102466
rect 45226 102418 45232 102426
rect 43378 102382 45232 102418
rect 45226 102374 45232 102382
rect 45284 102418 45290 102426
rect 45284 102382 45305 102418
rect 45284 102374 45290 102382
rect 45142 102334 45148 102343
rect 43378 102298 45148 102334
rect 45142 102291 45148 102298
rect 45200 102334 45206 102343
rect 45200 102298 45215 102334
rect 45200 102291 45206 102298
rect 45058 102250 45064 102258
rect 43378 102214 45064 102250
rect 45058 102206 45064 102214
rect 45116 102250 45122 102258
rect 45116 102214 45135 102250
rect 45116 102206 45122 102214
rect 44974 102166 44980 102173
rect 43378 102130 44980 102166
rect 44974 102121 44980 102130
rect 45032 102166 45038 102173
rect 45032 102130 45042 102166
rect 48330 102150 48410 102156
rect 45032 102121 45038 102130
rect 46906 102082 46912 102091
rect 43378 102046 46912 102082
rect 46906 102039 46912 102046
rect 46964 102082 46970 102091
rect 46964 102046 46974 102082
rect 48330 102064 48410 102070
rect 46964 102039 46970 102046
rect 46822 101998 46828 102007
rect 43378 101962 46828 101998
rect 46822 101955 46828 101962
rect 46880 101998 46886 102007
rect 46880 101962 46890 101998
rect 46880 101955 46886 101962
rect 46738 101914 46744 101922
rect 43378 101878 46744 101914
rect 46738 101870 46744 101878
rect 46796 101914 46802 101922
rect 46796 101878 46805 101914
rect 46796 101870 46802 101878
rect 46654 101830 46660 101838
rect 43378 101794 46660 101830
rect 46654 101786 46660 101794
rect 46712 101830 46718 101838
rect 46712 101794 46719 101830
rect 46712 101786 46718 101794
rect 46570 101746 46576 101755
rect 43378 101710 46576 101746
rect 46570 101703 46576 101710
rect 46628 101746 46634 101755
rect 46628 101710 46642 101746
rect 46628 101703 46634 101710
rect 46486 101662 46492 101672
rect 43378 101626 46492 101662
rect 46486 101620 46492 101626
rect 46544 101662 46550 101672
rect 46544 101626 46555 101662
rect 46544 101620 46550 101626
rect 48253 99786 48289 99791
rect 48230 99780 48310 99786
rect 48230 99694 48310 99700
rect 48149 97386 48185 97388
rect 48120 97380 48200 97386
rect 48120 97294 48200 97300
rect 47410 96720 47416 96728
rect 43404 96684 47416 96720
rect 47410 96676 47416 96684
rect 47468 96720 47474 96728
rect 47468 96684 47482 96720
rect 47468 96676 47474 96684
rect 47326 96636 47332 96644
rect 43404 96600 47332 96636
rect 47326 96592 47332 96600
rect 47384 96636 47390 96644
rect 47384 96600 47395 96636
rect 47384 96592 47390 96600
rect 47242 96552 47248 96561
rect 43404 96516 47248 96552
rect 47242 96509 47248 96516
rect 47300 96552 47306 96561
rect 47300 96516 47311 96552
rect 47300 96509 47306 96516
rect 47158 96468 47164 96477
rect 43404 96432 47164 96468
rect 47158 96425 47164 96432
rect 47216 96468 47222 96477
rect 47216 96432 47229 96468
rect 47216 96425 47222 96432
rect 47074 96384 47080 96391
rect 43404 96348 47080 96384
rect 47074 96339 47080 96348
rect 47132 96384 47138 96391
rect 47132 96348 47142 96384
rect 47132 96339 47138 96348
rect 46990 96300 46996 96310
rect 43404 96264 46996 96300
rect 46990 96258 46996 96264
rect 47048 96300 47054 96310
rect 47048 96264 47061 96300
rect 47048 96258 47054 96264
rect 46402 96216 46408 96226
rect 43404 96180 46408 96216
rect 46402 96174 46408 96180
rect 46460 96216 46466 96226
rect 46460 96180 46474 96216
rect 46460 96174 46466 96180
rect 46318 96132 46324 96141
rect 43404 96096 46324 96132
rect 46318 96089 46324 96096
rect 46376 96132 46382 96141
rect 46376 96096 46388 96132
rect 46376 96089 46382 96096
rect 46234 96048 46240 96058
rect 43404 96012 46240 96048
rect 46234 96006 46240 96012
rect 46292 96048 46298 96058
rect 46292 96012 46302 96048
rect 46292 96006 46298 96012
rect 46150 95964 46156 95972
rect 43404 95928 46156 95964
rect 46150 95920 46156 95928
rect 46208 95964 46214 95972
rect 46208 95928 46220 95964
rect 46208 95920 46214 95928
rect 46066 95880 46072 95892
rect 43404 95844 46072 95880
rect 46066 95840 46072 95844
rect 46124 95880 46130 95892
rect 46124 95844 46135 95880
rect 46124 95840 46130 95844
rect 45982 95796 45988 95804
rect 43404 95760 45988 95796
rect 45982 95752 45988 95760
rect 46040 95796 46046 95804
rect 46040 95760 46052 95796
rect 46040 95752 46046 95760
rect 48045 94986 48081 94994
rect 48014 94980 48094 94986
rect 48014 94894 48094 94900
rect 45898 90854 45904 90861
rect 43378 90818 45904 90854
rect 45898 90809 45904 90818
rect 45956 90854 45962 90861
rect 45956 90818 45968 90854
rect 45956 90809 45962 90818
rect 45814 90770 45820 90780
rect 43378 90734 45820 90770
rect 45814 90728 45820 90734
rect 45872 90770 45878 90780
rect 45872 90734 45884 90770
rect 45872 90728 45878 90734
rect 45730 90686 45736 90695
rect 43378 90650 45736 90686
rect 45730 90643 45736 90650
rect 45788 90686 45794 90695
rect 45788 90650 45807 90686
rect 45788 90643 45794 90650
rect 45646 90602 45652 90611
rect 43378 90566 45652 90602
rect 45646 90559 45652 90566
rect 45704 90602 45710 90611
rect 45704 90566 45718 90602
rect 45704 90559 45710 90566
rect 45562 90518 45568 90527
rect 43378 90482 45568 90518
rect 45562 90475 45568 90482
rect 45620 90475 45626 90527
rect 45478 90434 45484 90443
rect 43378 90398 45484 90434
rect 45478 90391 45484 90398
rect 45536 90434 45542 90443
rect 45536 90398 45551 90434
rect 45536 90391 45542 90398
rect 47494 90350 47500 90360
rect 43378 90314 47500 90350
rect 47494 90308 47500 90314
rect 47552 90350 47558 90360
rect 47552 90314 47564 90350
rect 47552 90308 47558 90314
rect 47914 90266 47920 90274
rect 43378 90230 47920 90266
rect 47914 90222 47920 90230
rect 47972 90222 47978 90274
rect 47830 90182 47836 90190
rect 43378 90146 47836 90182
rect 47830 90138 47836 90146
rect 47888 90138 47894 90190
rect 47746 90098 47752 90106
rect 43378 90062 47752 90098
rect 47746 90054 47752 90062
rect 47804 90054 47810 90106
rect 47662 90014 47668 90022
rect 43378 89978 47668 90014
rect 47662 89970 47668 89978
rect 47720 89970 47726 90022
rect 47578 89930 47584 89938
rect 43378 89894 47584 89930
rect 47578 89886 47584 89894
rect 47636 89886 47642 89938
rect 48045 89373 48081 94894
rect 47645 89337 48081 89373
rect 47645 85366 47681 89337
rect 48149 89269 48185 97294
rect 47145 85330 47681 85366
rect 47749 89233 48185 89269
rect 10142 84052 10148 84104
rect 10200 84092 10206 84104
rect 10200 84064 12817 84092
rect 10200 84052 10206 84064
rect 10254 83926 10260 83978
rect 10312 83966 10318 83978
rect 10312 83938 12800 83966
rect 10312 83926 10318 83938
rect 10366 83804 10372 83856
rect 10424 83844 10430 83856
rect 10424 83816 12817 83844
rect 10424 83804 10430 83816
rect 10478 83689 10484 83741
rect 10536 83729 10542 83741
rect 10536 83701 12810 83729
rect 10536 83689 10542 83701
rect 9918 78142 9924 78194
rect 9976 78182 9982 78194
rect 9976 78154 12826 78182
rect 9976 78142 9982 78154
rect 10030 78013 10036 78065
rect 10088 78053 10094 78065
rect 10088 78025 12793 78053
rect 10088 78013 10094 78025
rect 9694 77901 9700 77953
rect 9752 77941 9758 77953
rect 9752 77913 12813 77941
rect 9752 77901 9758 77913
rect 9806 77777 9812 77829
rect 9864 77817 9870 77829
rect 9864 77789 12783 77817
rect 9864 77777 9870 77789
rect 28883 77365 28889 77375
rect 28880 77329 28889 77365
rect 28883 77323 28889 77329
rect 28941 77365 28947 77375
rect 47145 77365 47181 85330
rect 47749 85262 47785 89233
rect 48253 89165 48289 99694
rect 28941 77329 47181 77365
rect 47249 85226 47785 85262
rect 47853 89129 48289 89165
rect 28941 77323 28947 77329
rect 28967 77281 28973 77291
rect 28964 77245 28973 77281
rect 28967 77239 28973 77245
rect 29025 77281 29031 77291
rect 47249 77281 47285 85226
rect 47853 85158 47889 89129
rect 48357 89061 48393 102064
rect 29025 77245 47285 77281
rect 47353 85122 47889 85158
rect 47957 89025 48393 89061
rect 29025 77239 29031 77245
rect 29051 77197 29057 77207
rect 29048 77161 29057 77197
rect 29051 77155 29057 77161
rect 29109 77197 29115 77207
rect 47353 77197 47389 85122
rect 47957 85054 47993 89025
rect 48461 88957 48497 104464
rect 286463 102999 286469 103061
rect 286531 102999 288103 103061
rect 286385 102768 288088 102775
rect 286383 102716 286389 102768
rect 286441 102716 288088 102768
rect 286385 102712 288088 102716
rect 508856 102554 508892 102561
rect 508830 102548 508910 102554
rect 508830 102462 508910 102468
rect 287308 101124 287314 101176
rect 287366 101168 287372 101176
rect 287366 101132 288057 101168
rect 287366 101124 287372 101132
rect 287224 101040 287230 101092
rect 287282 101084 287288 101092
rect 287282 101048 288057 101084
rect 287282 101040 287288 101048
rect 287727 100957 287733 101009
rect 287785 101000 287791 101009
rect 287785 100964 288059 101000
rect 287785 100957 287791 100964
rect 287811 100875 287817 100927
rect 287869 100916 287875 100927
rect 287869 100880 288059 100916
rect 287869 100875 287875 100880
rect 287055 100789 287061 100841
rect 287113 100832 287119 100841
rect 287113 100796 288063 100832
rect 287113 100789 287119 100796
rect 287139 100748 287145 100756
rect 287136 100712 287145 100748
rect 287139 100704 287145 100712
rect 287197 100748 287203 100756
rect 287197 100712 288063 100748
rect 287197 100704 287203 100712
rect 508762 100174 508798 100185
rect 508740 100168 508820 100174
rect 508740 100082 508820 100088
rect 508668 97758 508704 97770
rect 508642 97752 508722 97758
rect 508642 97666 508722 97672
rect 286887 93253 286893 93305
rect 286945 93298 286951 93305
rect 286945 93262 288070 93298
rect 286945 93253 286951 93262
rect 286970 93172 286977 93224
rect 287029 93214 287035 93224
rect 287029 93178 288070 93214
rect 287029 93172 287035 93178
rect 287474 93086 287480 93138
rect 287532 93130 287538 93138
rect 287532 93094 288062 93130
rect 287532 93086 287538 93094
rect 287392 93002 287398 93054
rect 287450 93046 287456 93054
rect 287450 93010 288062 93046
rect 287450 93002 287456 93010
rect 287559 92917 287565 92969
rect 287617 92962 287623 92969
rect 287617 92926 288065 92962
rect 287617 92917 287623 92926
rect 287643 92878 287649 92888
rect 287642 92842 287649 92878
rect 287643 92836 287649 92842
rect 287701 92878 287707 92888
rect 287701 92842 288065 92878
rect 287701 92836 287707 92842
rect 48550 92569 48602 92575
rect 48550 92511 48602 92517
rect 48558 90806 48594 92511
rect 434140 90895 435650 90933
rect 388877 90856 390307 90889
rect 48558 90770 48717 90806
rect 48532 90180 48612 90186
rect 48532 90094 48612 90100
rect 29109 77161 47389 77197
rect 47457 85018 47993 85054
rect 48061 88921 48497 88957
rect 48558 90078 48595 90094
rect 29109 77155 29115 77161
rect 29135 77113 29141 77123
rect 29132 77077 29141 77113
rect 29135 77071 29141 77077
rect 29193 77113 29199 77123
rect 47457 77113 47493 85018
rect 48061 84950 48097 88921
rect 48558 88596 48594 90078
rect 48477 88560 48594 88596
rect 48365 87746 48417 87752
rect 48365 87688 48417 87694
rect 48269 85376 48305 85393
rect 48261 85370 48313 85376
rect 48261 85312 48313 85318
rect 29193 77077 47493 77113
rect 47561 84914 48097 84950
rect 29193 77071 29199 77077
rect 29219 77029 29225 77039
rect 29216 76993 29225 77029
rect 29219 76987 29225 76993
rect 29277 77029 29283 77039
rect 47561 77029 47597 84914
rect 48165 82972 48201 82978
rect 48157 82966 48213 82972
rect 48157 82904 48213 82910
rect 29277 76993 47597 77029
rect 29277 76987 29283 76993
rect 29303 76945 29309 76955
rect 29300 76909 29309 76945
rect 29303 76903 29309 76909
rect 29361 76945 29367 76955
rect 48165 76945 48201 82904
rect 29361 76909 48201 76945
rect 29361 76903 29367 76909
rect 29387 76861 29393 76871
rect 29384 76825 29393 76861
rect 29387 76819 29393 76825
rect 29445 76861 29451 76871
rect 48269 76861 48305 85312
rect 29445 76825 48305 76861
rect 29445 76819 29451 76825
rect 29471 76777 29477 76787
rect 29468 76741 29477 76777
rect 29471 76735 29477 76741
rect 29529 76777 29535 76787
rect 48373 76777 48409 87688
rect 29529 76741 48409 76777
rect 29529 76735 29535 76741
rect 29555 76693 29561 76703
rect 29552 76657 29561 76693
rect 29555 76651 29561 76657
rect 29613 76693 29619 76703
rect 48477 76693 48513 88560
rect 48681 88364 48717 90770
rect 388877 90725 388908 90856
rect 390258 90725 390307 90856
rect 434140 90780 434187 90895
rect 435612 90780 435650 90895
rect 434140 90741 435650 90780
rect 388877 90694 390307 90725
rect 198816 90609 200403 90635
rect 198816 90469 198858 90609
rect 200372 90469 200403 90609
rect 198816 90451 200403 90469
rect 154532 90355 156082 90383
rect 154532 90232 154585 90355
rect 156040 90232 156082 90355
rect 154532 90196 156082 90232
rect 434430 90110 435108 90146
rect 389468 90071 390701 90107
rect 196216 89834 196222 89886
rect 196274 89878 196280 89886
rect 196274 89842 199868 89878
rect 196274 89834 196280 89842
rect 158300 89643 158352 89649
rect 155131 89599 158300 89635
rect 158300 89585 158352 89591
rect 388959 89308 390389 89349
rect 388959 89177 388995 89308
rect 390345 89177 390389 89308
rect 388959 89154 390389 89177
rect 198818 89070 200387 89093
rect 198818 88930 198845 89070
rect 200359 88930 200387 89070
rect 198818 88915 200387 88930
rect 154634 88824 156048 88857
rect 154634 88696 154673 88824
rect 156003 88696 156048 88824
rect 154634 88671 156048 88696
rect 29613 76657 48513 76693
rect 48581 88328 48717 88364
rect 29613 76651 29619 76657
rect 29639 76609 29645 76619
rect 29636 76573 29645 76609
rect 29639 76567 29645 76573
rect 29697 76609 29703 76619
rect 48581 76609 48617 88328
rect 286630 86946 286636 87006
rect 286696 86946 288050 87006
rect 286562 86702 288089 86710
rect 286551 86650 286557 86702
rect 286609 86650 288089 86702
rect 286562 86649 288089 86650
rect 286804 85048 286810 85100
rect 286862 85092 286868 85100
rect 286862 85056 288077 85092
rect 286862 85048 286868 85056
rect 286719 84964 286725 85016
rect 286777 85008 286783 85016
rect 286777 84972 288077 85008
rect 286777 84964 286783 84972
rect 287140 84880 287146 84932
rect 287198 84924 287204 84932
rect 287198 84888 288077 84924
rect 287198 84880 287204 84888
rect 287056 84796 287062 84848
rect 287114 84840 287120 84848
rect 287114 84804 288077 84840
rect 287114 84796 287120 84804
rect 289599 84712 289605 84764
rect 289657 84712 289663 84764
rect 289683 84627 289689 84679
rect 289741 84627 289747 84679
rect 287979 83284 287985 83336
rect 288037 83329 288043 83336
rect 289011 83329 289017 83338
rect 288037 83293 289017 83329
rect 288037 83284 288043 83293
rect 289011 83286 289017 83293
rect 289069 83286 289075 83338
rect 287895 83200 287901 83252
rect 287953 83245 287959 83252
rect 288927 83245 288933 83254
rect 287953 83209 288933 83245
rect 287953 83200 287959 83209
rect 288927 83202 288933 83209
rect 288985 83202 288991 83254
rect 287811 83116 287817 83168
rect 287869 83161 287875 83168
rect 288843 83161 288849 83170
rect 287869 83125 288849 83161
rect 287869 83116 287875 83125
rect 288843 83118 288849 83125
rect 288901 83118 288907 83170
rect 287727 83032 287733 83084
rect 287785 83077 287791 83084
rect 288759 83077 288765 83086
rect 287785 83041 288765 83077
rect 287785 83032 287791 83041
rect 288759 83034 288765 83041
rect 288817 83034 288823 83086
rect 287307 82949 287313 83001
rect 287365 82993 287371 83001
rect 288339 82993 288345 83000
rect 287365 82957 288345 82993
rect 287365 82949 287371 82957
rect 288339 82948 288345 82957
rect 288397 82948 288403 83000
rect 287223 82865 287229 82917
rect 287281 82909 287287 82917
rect 288255 82909 288261 82916
rect 287281 82873 288261 82909
rect 287281 82865 287287 82873
rect 288255 82864 288261 82873
rect 288313 82864 288319 82916
rect 286971 82782 286977 82834
rect 287029 82825 287035 82834
rect 288171 82825 288177 82832
rect 287029 82789 288177 82825
rect 287029 82782 287035 82789
rect 288171 82780 288177 82789
rect 288229 82780 288235 82832
rect 286887 82698 286893 82750
rect 286945 82741 286951 82750
rect 288087 82741 288093 82748
rect 286945 82705 288093 82741
rect 286945 82698 286951 82705
rect 288087 82696 288093 82705
rect 288145 82696 288151 82748
rect 48747 81227 49085 81245
rect 48747 80907 48765 81227
rect 49066 80907 49085 81227
rect 48747 80887 49085 80907
rect 48747 79997 49083 80015
rect 48747 79677 48765 79997
rect 49066 79677 49083 79997
rect 48747 79660 49083 79677
rect 163163 78030 163169 78038
rect 29697 76573 48617 76609
rect 93241 77994 163169 78030
rect 29697 76567 29703 76573
rect 29723 76525 29729 76535
rect 29720 76489 29729 76525
rect 29723 76483 29729 76489
rect 29781 76525 29787 76535
rect 93241 76525 93277 77994
rect 163163 77986 163169 77994
rect 163221 77986 163227 78038
rect 158294 77946 158300 77955
rect 29781 76489 93277 76525
rect 93325 77910 158300 77946
rect 29781 76483 29787 76489
rect 29807 76441 29813 76451
rect 29804 76405 29813 76441
rect 29807 76399 29813 76405
rect 29865 76441 29871 76451
rect 93325 76441 93361 77910
rect 158294 77903 158300 77910
rect 158352 77946 158358 77955
rect 158352 77910 158366 77946
rect 158352 77903 158358 77910
rect 94224 77827 94230 77835
rect 94220 77791 94230 77827
rect 94224 77783 94230 77791
rect 94282 77827 94288 77835
rect 163349 77827 163407 81173
rect 94282 77791 163407 77827
rect 94282 77783 94288 77791
rect 94308 77743 94314 77751
rect 94304 77707 94314 77743
rect 94308 77699 94314 77707
rect 94366 77743 94372 77751
rect 164977 77743 165035 81148
rect 94366 77707 165035 77743
rect 94366 77699 94372 77707
rect 94392 77659 94398 77667
rect 94388 77623 94398 77659
rect 94392 77615 94398 77623
rect 94450 77659 94456 77667
rect 166605 77659 166663 81163
rect 94450 77623 166663 77659
rect 94450 77615 94456 77623
rect 94476 77575 94482 77583
rect 94472 77539 94482 77575
rect 94476 77531 94482 77539
rect 94534 77575 94540 77583
rect 168233 77575 168291 81148
rect 94534 77539 168291 77575
rect 94534 77531 94540 77539
rect 94560 77491 94566 77499
rect 94556 77455 94566 77491
rect 94560 77447 94566 77455
rect 94618 77491 94624 77499
rect 169861 77491 169919 81179
rect 94618 77455 169919 77491
rect 94618 77447 94624 77455
rect 94644 77407 94650 77415
rect 94640 77371 94650 77407
rect 94644 77363 94650 77371
rect 94702 77407 94708 77415
rect 171489 77407 171547 81185
rect 94702 77371 171547 77407
rect 94702 77363 94708 77371
rect 94728 77323 94734 77331
rect 94724 77287 94734 77323
rect 94728 77279 94734 77287
rect 94786 77323 94792 77331
rect 173117 77323 173175 81148
rect 94786 77287 173175 77323
rect 94786 77279 94792 77287
rect 94812 77239 94818 77247
rect 94808 77203 94818 77239
rect 94812 77195 94818 77203
rect 94870 77239 94876 77247
rect 174745 77239 174803 81148
rect 94870 77203 174803 77239
rect 94870 77195 94876 77203
rect 94896 77155 94902 77163
rect 94892 77119 94902 77155
rect 94896 77111 94902 77119
rect 94954 77155 94960 77163
rect 179817 77155 179875 81130
rect 94954 77119 179875 77155
rect 94954 77111 94960 77119
rect 94980 77071 94986 77079
rect 94976 77035 94986 77071
rect 94980 77027 94986 77035
rect 95038 77071 95044 77079
rect 181445 77071 181503 81130
rect 95038 77035 181503 77071
rect 95038 77027 95044 77035
rect 95064 76987 95070 76995
rect 95060 76951 95070 76987
rect 95064 76943 95070 76951
rect 95122 76987 95128 76995
rect 183073 76987 183131 81130
rect 95122 76951 183131 76987
rect 95122 76943 95128 76951
rect 95148 76903 95154 76911
rect 95144 76867 95154 76903
rect 95148 76859 95154 76867
rect 95206 76903 95212 76911
rect 184701 76903 184759 81137
rect 95206 76867 184759 76903
rect 95206 76859 95212 76867
rect 95232 76819 95238 76827
rect 95228 76783 95238 76819
rect 95232 76775 95238 76783
rect 95290 76819 95296 76827
rect 186329 76819 186387 81159
rect 95290 76783 186387 76819
rect 95290 76775 95296 76783
rect 95316 76735 95322 76743
rect 95312 76699 95322 76735
rect 95316 76691 95322 76699
rect 95374 76735 95380 76743
rect 187957 76735 188015 81158
rect 95374 76699 188015 76735
rect 95374 76691 95380 76699
rect 95400 76651 95406 76659
rect 95396 76615 95406 76651
rect 95400 76607 95406 76615
rect 95458 76651 95464 76659
rect 189585 76651 189643 81138
rect 95458 76615 189643 76651
rect 95458 76607 95464 76615
rect 95484 76567 95490 76575
rect 95480 76531 95490 76567
rect 95484 76523 95490 76531
rect 95542 76567 95548 76575
rect 191213 76567 191271 81142
rect 390665 79049 390701 90071
rect 434430 84381 434466 90110
rect 434605 89395 435575 89397
rect 434605 89367 436007 89395
rect 434605 89231 434639 89367
rect 435961 89231 436007 89367
rect 434605 89197 436007 89231
rect 434430 84345 507603 84381
rect 431330 84243 507481 84279
rect 397727 79166 397785 80718
rect 399355 79250 399413 80700
rect 400983 79334 401041 80696
rect 402611 79418 402669 80696
rect 404239 79502 404297 80696
rect 405867 79586 405925 80696
rect 407495 79670 407553 80696
rect 409123 79754 409181 80696
rect 413895 79838 413953 80636
rect 415523 79922 415581 80636
rect 417151 80006 417209 80636
rect 418779 80090 418837 80636
rect 420407 80174 420465 80636
rect 422035 80258 422093 80636
rect 423663 80342 423721 80636
rect 425291 80426 425349 80685
rect 431330 80426 431366 84243
rect 425291 80390 431366 80426
rect 431414 84159 507397 84195
rect 431414 80342 431450 84159
rect 423663 80306 431450 80342
rect 431498 84075 507313 84111
rect 431498 80258 431534 84075
rect 422035 80222 431534 80258
rect 431582 83991 507229 84027
rect 431582 80174 431618 83991
rect 420407 80138 431618 80174
rect 431666 83907 507145 83943
rect 431666 80090 431702 83907
rect 418779 80054 431702 80090
rect 431750 83823 507061 83859
rect 431750 80006 431786 83823
rect 417151 79970 431786 80006
rect 431834 83739 506977 83775
rect 431834 79922 431870 83739
rect 415523 79886 431870 79922
rect 431918 83655 506893 83691
rect 431918 79838 431954 83655
rect 413895 79802 431954 79838
rect 432002 83571 506809 83607
rect 432002 79754 432038 83571
rect 409123 79718 432038 79754
rect 432086 83487 506725 83523
rect 432086 79670 432122 83487
rect 407495 79634 432122 79670
rect 432170 83403 506641 83439
rect 432170 79586 432206 83403
rect 405867 79550 432206 79586
rect 432254 83319 506557 83355
rect 432254 79502 432290 83319
rect 404239 79466 432290 79502
rect 432338 83235 506473 83271
rect 432338 79418 432374 83235
rect 402611 79382 432374 79418
rect 432422 83151 506389 83187
rect 432422 79334 432458 83151
rect 400983 79298 432458 79334
rect 432506 83067 506305 83103
rect 432506 79250 432542 83067
rect 399355 79214 432542 79250
rect 432590 82983 506221 83019
rect 432590 79166 432626 82983
rect 397727 79130 432626 79166
rect 432681 82880 506130 82916
rect 432681 79049 432717 82880
rect 390665 79013 432717 79049
rect 506094 78581 506130 82880
rect 506185 78672 506221 82983
rect 506269 78756 506305 83067
rect 506353 78840 506389 83151
rect 506437 78924 506473 83235
rect 506521 79008 506557 83319
rect 506605 79092 506641 83403
rect 506689 79176 506725 83487
rect 506773 79260 506809 83571
rect 506857 79344 506893 83655
rect 506941 79428 506977 83739
rect 507025 79512 507061 83823
rect 507109 79596 507145 83907
rect 507193 79680 507229 83991
rect 507277 79764 507313 84075
rect 507361 79848 507397 84159
rect 507445 79932 507481 84243
rect 507567 80037 507603 84345
rect 507567 80001 508292 80037
rect 507532 79932 507538 79940
rect 507445 79896 507538 79932
rect 507532 79888 507538 79896
rect 507590 79888 507596 79940
rect 507616 79848 507622 79857
rect 507361 79812 507622 79848
rect 507616 79805 507622 79812
rect 507674 79848 507680 79857
rect 507674 79812 507682 79848
rect 507674 79805 507680 79812
rect 507701 79764 507707 79773
rect 507277 79728 507707 79764
rect 507701 79721 507707 79728
rect 507759 79764 507765 79773
rect 507759 79728 507766 79764
rect 507759 79721 507765 79728
rect 507785 79680 507791 79688
rect 507193 79644 507791 79680
rect 507785 79636 507791 79644
rect 507843 79680 507849 79688
rect 507843 79644 507850 79680
rect 507843 79636 507849 79644
rect 507869 79596 507875 79604
rect 507109 79560 507875 79596
rect 507869 79552 507875 79560
rect 507927 79596 507933 79604
rect 507927 79560 507934 79596
rect 507927 79552 507933 79560
rect 507953 79512 507959 79521
rect 507025 79476 507959 79512
rect 507953 79469 507959 79476
rect 508011 79512 508017 79521
rect 508011 79476 508018 79512
rect 508011 79469 508017 79476
rect 508037 79428 508043 79435
rect 506941 79392 508043 79428
rect 508037 79383 508043 79392
rect 508095 79428 508101 79435
rect 508095 79392 508102 79428
rect 508095 79383 508101 79392
rect 508121 79344 508127 79352
rect 506857 79308 508127 79344
rect 508121 79300 508127 79308
rect 508179 79344 508185 79352
rect 508179 79308 508186 79344
rect 508179 79300 508185 79308
rect 507448 79260 507454 79269
rect 506765 79224 507454 79260
rect 507448 79217 507454 79224
rect 507506 79260 507512 79269
rect 507506 79224 507523 79260
rect 507506 79217 507512 79224
rect 507364 79176 507370 79185
rect 506689 79140 507370 79176
rect 507364 79133 507370 79140
rect 507422 79176 507428 79185
rect 507422 79140 507439 79176
rect 507422 79133 507428 79140
rect 507280 79092 507286 79101
rect 506605 79056 507286 79092
rect 507280 79049 507286 79056
rect 507338 79092 507344 79101
rect 507338 79056 507355 79092
rect 507338 79049 507344 79056
rect 507196 79008 507202 79017
rect 506521 78972 507202 79008
rect 507196 78965 507202 78972
rect 507254 79008 507260 79017
rect 507254 78972 507271 79008
rect 507254 78965 507260 78972
rect 507112 78924 507118 78933
rect 506437 78888 507118 78924
rect 507112 78881 507118 78888
rect 507170 78924 507176 78933
rect 507170 78888 507187 78924
rect 507170 78881 507176 78888
rect 507028 78840 507034 78849
rect 506353 78804 507034 78840
rect 507028 78797 507034 78804
rect 507086 78840 507092 78849
rect 507086 78804 507103 78840
rect 507086 78797 507092 78804
rect 506944 78756 506950 78765
rect 506269 78720 506950 78756
rect 506944 78713 506950 78720
rect 507002 78756 507008 78765
rect 507002 78720 507019 78756
rect 507002 78713 507008 78720
rect 506860 78672 506866 78681
rect 506185 78636 506866 78672
rect 506860 78629 506866 78636
rect 506918 78672 506924 78681
rect 508256 78677 508292 80001
rect 508668 79053 508704 97666
rect 508762 79147 508798 100082
rect 508856 79241 508892 102462
rect 508950 79335 508986 104860
rect 509044 79429 509080 107268
rect 509514 95368 509550 95371
rect 509485 95362 509565 95368
rect 509485 95276 509565 95282
rect 509420 92978 509456 92980
rect 509398 92972 509478 92978
rect 509398 92886 509478 92892
rect 509326 90568 509362 90571
rect 509303 90562 509383 90568
rect 509303 90476 509383 90482
rect 509238 88177 509274 88181
rect 509230 88171 509282 88177
rect 509230 88113 509282 88119
rect 509155 85760 509191 85788
rect 509147 85754 509199 85760
rect 509147 85696 509199 85702
rect 509155 79534 509191 85696
rect 509238 79618 509274 88113
rect 509326 79711 509362 90476
rect 509420 79805 509456 92886
rect 509514 79899 509550 95276
rect 568818 88974 568824 88986
rect 568584 88946 568824 88974
rect 568818 88934 568824 88946
rect 568876 88934 568882 88986
rect 568930 88860 568936 88872
rect 568614 88832 568936 88860
rect 568930 88820 568936 88832
rect 568988 88820 568994 88872
rect 569042 88740 569048 88752
rect 568598 88712 569048 88740
rect 569042 88700 569048 88712
rect 569100 88700 569106 88752
rect 569154 88606 569160 88618
rect 568604 88578 569160 88606
rect 569154 88566 569160 88578
rect 569212 88566 569218 88618
rect 509741 83844 510994 83859
rect 509741 83681 509759 83844
rect 510920 83681 510994 83844
rect 509741 83662 510994 83681
rect 569266 83062 569272 83074
rect 568604 83034 569272 83062
rect 569266 83022 569272 83034
rect 569324 83022 569330 83074
rect 569378 82944 569384 82956
rect 568574 82916 569384 82944
rect 569378 82904 569384 82916
rect 569436 82904 569442 82956
rect 569490 82824 569496 82836
rect 568598 82796 569496 82824
rect 569490 82784 569496 82796
rect 569548 82784 569554 82836
rect 509747 82704 510995 82720
rect 569602 82710 569608 82722
rect 509747 82541 509771 82704
rect 510932 82541 510995 82704
rect 568568 82682 569608 82710
rect 569602 82670 569608 82682
rect 569660 82670 569666 82722
rect 509747 82520 510995 82541
rect 509514 79863 511670 79899
rect 509420 79769 511576 79805
rect 509326 79675 511482 79711
rect 509238 79582 511388 79618
rect 509155 79498 511294 79534
rect 509044 79393 511200 79429
rect 508950 79299 511106 79335
rect 508856 79205 511012 79241
rect 508762 79111 510918 79147
rect 508668 79017 510824 79053
rect 506918 78636 506935 78672
rect 508256 78641 510646 78677
rect 506918 78629 506924 78636
rect 506094 78545 510562 78581
rect 510396 78446 510402 78454
rect 398166 78410 510402 78446
rect 376242 78362 376248 78376
rect 376227 78326 376248 78362
rect 376242 78324 376248 78326
rect 376300 78362 376306 78376
rect 398166 78362 398202 78410
rect 510396 78402 510402 78410
rect 510454 78446 510460 78454
rect 510454 78410 510462 78446
rect 510454 78402 510460 78410
rect 510312 78362 510318 78370
rect 376300 78326 398202 78362
rect 398340 78326 510318 78362
rect 376300 78324 376306 78326
rect 380660 78278 380666 78279
rect 380649 78242 380666 78278
rect 380660 78227 380666 78242
rect 380718 78278 380724 78279
rect 398340 78278 398376 78326
rect 510312 78318 510318 78326
rect 510370 78362 510376 78370
rect 510370 78326 510378 78362
rect 510370 78318 510376 78326
rect 458764 78278 458770 78282
rect 380718 78242 398376 78278
rect 458754 78242 458770 78278
rect 380718 78227 380724 78242
rect 458764 78230 458770 78242
rect 458822 78278 458828 78282
rect 510228 78278 510234 78286
rect 458822 78242 510234 78278
rect 458822 78230 458828 78242
rect 510228 78234 510234 78242
rect 510286 78278 510292 78286
rect 510286 78242 510294 78278
rect 510286 78234 510292 78242
rect 385194 78194 385200 78197
rect 385182 78158 385200 78194
rect 385194 78145 385200 78158
rect 385252 78194 385258 78197
rect 510144 78194 510150 78202
rect 385252 78158 510150 78194
rect 385252 78145 385258 78158
rect 510144 78150 510150 78158
rect 510202 78194 510208 78202
rect 510202 78158 510210 78194
rect 510202 78150 510208 78158
rect 482236 78110 482242 78118
rect 482223 78074 482242 78110
rect 482236 78066 482242 78074
rect 482294 78110 482300 78118
rect 510060 78110 510066 78118
rect 482294 78074 510066 78110
rect 482294 78066 482300 78074
rect 510060 78066 510066 78074
rect 510118 78110 510124 78118
rect 510118 78074 510126 78110
rect 510118 78066 510124 78074
rect 191486 78038 191538 78044
rect 196216 78030 196222 78038
rect 191538 77994 196222 78030
rect 196216 77986 196222 77994
rect 196274 77986 196280 78038
rect 445184 78026 445190 78040
rect 445176 77990 445190 78026
rect 445184 77988 445190 77990
rect 445242 78026 445248 78040
rect 509976 78026 509982 78034
rect 445242 77990 509982 78026
rect 445242 77988 445248 77990
rect 191486 77980 191538 77986
rect 509976 77982 509982 77990
rect 510034 78026 510040 78034
rect 510034 77990 510042 78026
rect 510034 77982 510040 77990
rect 440450 77942 440456 77948
rect 440444 77906 440456 77942
rect 440450 77896 440456 77906
rect 440508 77942 440514 77948
rect 509892 77942 509898 77950
rect 440508 77906 509898 77942
rect 440508 77896 440514 77906
rect 509892 77898 509898 77906
rect 509950 77942 509956 77950
rect 509950 77906 509958 77942
rect 509950 77898 509956 77906
rect 454378 77858 454384 77864
rect 454366 77822 454384 77858
rect 454378 77812 454384 77822
rect 454436 77858 454442 77864
rect 509808 77858 509814 77866
rect 454436 77822 509814 77858
rect 454436 77812 454442 77822
rect 509808 77814 509814 77822
rect 509866 77858 509872 77866
rect 509866 77822 509874 77858
rect 509866 77814 509872 77822
rect 435832 77774 435838 77776
rect 435820 77738 435838 77774
rect 435832 77724 435838 77738
rect 435890 77774 435896 77776
rect 509724 77774 509730 77782
rect 435890 77738 509730 77774
rect 435890 77724 435896 77738
rect 509724 77730 509730 77738
rect 509782 77774 509788 77782
rect 509782 77738 509790 77774
rect 509782 77730 509788 77738
rect 477520 77690 477526 77696
rect 477506 77654 477526 77690
rect 477520 77644 477526 77654
rect 477578 77690 477584 77696
rect 509640 77690 509646 77698
rect 477578 77654 509646 77690
rect 477578 77644 477584 77654
rect 509640 77646 509646 77654
rect 509698 77690 509704 77698
rect 509698 77654 509706 77690
rect 509698 77646 509704 77654
rect 463580 77606 463586 77616
rect 463568 77570 463586 77606
rect 463580 77564 463586 77570
rect 463638 77606 463644 77616
rect 509556 77606 509562 77614
rect 463638 77570 509562 77606
rect 463638 77564 463644 77570
rect 509556 77562 509562 77570
rect 509614 77606 509620 77614
rect 509614 77570 509622 77606
rect 509614 77562 509620 77570
rect 486852 77522 486858 77532
rect 486844 77486 486858 77522
rect 486852 77480 486858 77486
rect 486910 77522 486916 77532
rect 509472 77522 509478 77530
rect 486910 77486 509478 77522
rect 486910 77480 486916 77486
rect 509472 77478 509478 77486
rect 509530 77522 509536 77530
rect 509530 77486 509538 77522
rect 509530 77478 509536 77486
rect 468226 77438 468232 77444
rect 468218 77402 468232 77438
rect 468226 77392 468232 77402
rect 468284 77438 468290 77444
rect 509388 77438 509394 77446
rect 468284 77402 509394 77438
rect 468284 77392 468290 77402
rect 509388 77394 509394 77402
rect 509446 77438 509452 77446
rect 509446 77402 509454 77438
rect 509446 77394 509452 77402
rect 491468 77354 491474 77364
rect 491460 77318 491474 77354
rect 491468 77312 491474 77318
rect 491526 77354 491532 77364
rect 509304 77354 509310 77362
rect 491526 77318 509310 77354
rect 491526 77312 491532 77318
rect 509304 77310 509310 77318
rect 509362 77354 509368 77362
rect 509362 77318 509370 77354
rect 509362 77310 509368 77318
rect 510526 77271 510562 78545
rect 510610 77367 510646 78641
rect 510788 77547 510824 79017
rect 510882 77631 510918 79111
rect 510976 77715 511012 79205
rect 511070 77799 511106 79299
rect 511164 77883 511200 79393
rect 511258 77967 511294 79498
rect 511352 78051 511388 79582
rect 511446 78135 511482 79675
rect 511540 78219 511576 79769
rect 511634 78303 511670 79863
rect 528464 78303 528470 78310
rect 511634 78267 528470 78303
rect 528464 78258 528470 78267
rect 528522 78303 528528 78310
rect 528522 78267 528534 78303
rect 528522 78258 528528 78267
rect 528380 78219 528386 78226
rect 511540 78183 528386 78219
rect 528380 78174 528386 78183
rect 528438 78219 528444 78226
rect 528438 78183 528450 78219
rect 528438 78174 528444 78183
rect 528296 78135 528302 78142
rect 511446 78099 528302 78135
rect 528296 78090 528302 78099
rect 528354 78135 528360 78142
rect 528354 78099 528366 78135
rect 528354 78090 528360 78099
rect 528212 78051 528218 78058
rect 511352 78015 528218 78051
rect 528212 78006 528218 78015
rect 528270 78051 528276 78058
rect 528270 78015 528282 78051
rect 528270 78006 528276 78015
rect 528128 77967 528134 77974
rect 511258 77931 528134 77967
rect 528128 77922 528134 77931
rect 528186 77967 528192 77974
rect 528186 77931 528198 77967
rect 528186 77922 528192 77931
rect 528044 77883 528050 77890
rect 511164 77847 528050 77883
rect 528044 77838 528050 77847
rect 528102 77883 528108 77890
rect 528102 77847 528114 77883
rect 528102 77838 528108 77847
rect 527960 77799 527966 77806
rect 511070 77763 527966 77799
rect 527960 77754 527966 77763
rect 528018 77799 528024 77806
rect 528018 77763 528030 77799
rect 528018 77754 528024 77763
rect 527876 77715 527882 77722
rect 510976 77679 527882 77715
rect 527876 77670 527882 77679
rect 527934 77715 527940 77722
rect 527934 77679 527946 77715
rect 527934 77670 527940 77679
rect 527792 77631 527798 77638
rect 510882 77595 527798 77631
rect 527792 77586 527798 77595
rect 527850 77631 527856 77638
rect 527850 77595 527862 77631
rect 527850 77586 527856 77595
rect 527708 77547 527714 77554
rect 510788 77511 527714 77547
rect 527708 77502 527714 77511
rect 527766 77547 527772 77554
rect 527766 77511 527778 77547
rect 527766 77502 527772 77511
rect 528632 77367 528638 77375
rect 510610 77331 528638 77367
rect 528632 77323 528638 77331
rect 528690 77323 528696 77375
rect 528551 77271 528557 77279
rect 510526 77235 528557 77271
rect 289431 77178 289437 77230
rect 289489 77178 289495 77230
rect 528551 77227 528557 77235
rect 528609 77227 528615 77279
rect 527408 77184 527414 77192
rect 367570 77148 527414 77184
rect 289515 77094 289521 77146
rect 289573 77094 289579 77146
rect 286972 77010 286978 77062
rect 287030 77054 287036 77062
rect 287030 77018 288061 77054
rect 287030 77010 287036 77018
rect 286888 76926 286894 76978
rect 286946 76970 286952 76978
rect 286946 76934 288061 76970
rect 286946 76926 286952 76934
rect 287306 76842 287312 76894
rect 287364 76886 287370 76894
rect 287364 76850 288062 76886
rect 287364 76842 287370 76850
rect 287223 76758 287229 76810
rect 287281 76802 287287 76810
rect 287281 76766 288062 76802
rect 287281 76758 287287 76766
rect 95542 76531 191271 76567
rect 95542 76523 95548 76531
rect 29865 76405 93361 76441
rect 29865 76399 29871 76405
rect 34590 76025 34596 76077
rect 34648 76069 34654 76077
rect 231372 76069 231378 76076
rect 34648 76033 231378 76069
rect 34648 76025 34654 76033
rect 231372 76024 231378 76033
rect 231430 76069 231436 76076
rect 231430 76033 231443 76069
rect 231430 76024 231436 76033
rect 34674 75985 34680 75993
rect 34670 75949 34680 75985
rect 34674 75941 34680 75949
rect 34732 75985 34738 75993
rect 199058 75985 199064 75998
rect 34732 75949 199064 75985
rect 34732 75941 34738 75949
rect 199058 75946 199064 75949
rect 199116 75985 199122 75998
rect 199116 75949 199124 75985
rect 199116 75946 199122 75949
rect 34758 75901 34764 75909
rect 34754 75865 34764 75901
rect 34758 75857 34764 75865
rect 34816 75901 34822 75909
rect 219886 75901 219892 75912
rect 34816 75865 219892 75901
rect 34816 75857 34822 75865
rect 219886 75860 219892 75865
rect 219944 75901 219950 75912
rect 219944 75865 219963 75901
rect 219944 75860 219950 75865
rect 34842 75817 34848 75825
rect 34838 75781 34848 75817
rect 34842 75773 34848 75781
rect 34900 75817 34906 75825
rect 203476 75817 203482 75831
rect 34900 75781 203482 75817
rect 34900 75773 34906 75781
rect 203476 75779 203482 75781
rect 203534 75817 203540 75831
rect 203534 75781 203551 75817
rect 203534 75779 203540 75781
rect 34926 75733 34932 75741
rect 34922 75697 34932 75733
rect 34926 75689 34932 75697
rect 34984 75733 34990 75741
rect 208010 75733 208016 75743
rect 34984 75697 208016 75733
rect 34984 75689 34990 75697
rect 208010 75691 208016 75697
rect 208068 75733 208074 75743
rect 208068 75697 208098 75733
rect 208068 75691 208074 75697
rect 35010 75649 35016 75657
rect 35006 75613 35016 75649
rect 35010 75605 35016 75613
rect 35068 75649 35074 75657
rect 235888 75649 235894 75660
rect 35068 75613 235894 75649
rect 35068 75605 35074 75613
rect 235888 75608 235894 75613
rect 235946 75649 235952 75660
rect 235946 75613 235965 75649
rect 235946 75608 235952 75613
rect 35094 75565 35100 75573
rect 35090 75529 35100 75565
rect 35094 75521 35100 75529
rect 35152 75565 35158 75573
rect 152448 75565 152454 75580
rect 35152 75529 152454 75565
rect 35152 75521 35158 75529
rect 152448 75528 152454 75529
rect 152506 75565 152512 75580
rect 152506 75529 152518 75565
rect 152506 75528 152512 75529
rect 35178 75481 35184 75489
rect 35174 75445 35184 75481
rect 35178 75437 35184 75445
rect 35236 75481 35242 75489
rect 224402 75481 224408 75490
rect 35236 75445 224408 75481
rect 35236 75437 35242 75445
rect 224402 75438 224408 75445
rect 224460 75481 224466 75490
rect 224460 75445 224490 75481
rect 224460 75438 224466 75445
rect 35262 75397 35268 75405
rect 35258 75361 35268 75397
rect 35262 75353 35268 75361
rect 35320 75397 35326 75405
rect 147914 75397 147920 75408
rect 35320 75361 147920 75397
rect 35320 75353 35326 75361
rect 147914 75356 147920 75361
rect 147972 75397 147978 75408
rect 147972 75361 148001 75397
rect 147972 75356 147978 75361
rect 147914 75351 147978 75356
rect 35346 75313 35352 75321
rect 35342 75277 35352 75313
rect 35346 75269 35352 75277
rect 35404 75313 35410 75321
rect 143496 75313 143502 75321
rect 35404 75277 143502 75313
rect 35404 75269 35410 75277
rect 143496 75269 143502 75277
rect 143554 75313 143560 75321
rect 143554 75277 143580 75313
rect 143554 75269 143560 75277
rect 35430 75229 35436 75237
rect 35426 75193 35436 75229
rect 35430 75185 35436 75193
rect 35488 75229 35494 75237
rect 240404 75229 240410 75235
rect 35488 75193 240410 75229
rect 35488 75185 35494 75193
rect 240404 75183 240410 75193
rect 240462 75229 240468 75235
rect 240462 75193 240484 75229
rect 240462 75183 240468 75193
rect 35514 75145 35520 75153
rect 35510 75109 35520 75145
rect 35514 75101 35520 75109
rect 35572 75145 35578 75153
rect 215370 75145 215376 75152
rect 35572 75109 215376 75145
rect 35572 75101 35578 75109
rect 215370 75100 215376 75109
rect 215428 75145 215434 75152
rect 215428 75109 215436 75145
rect 367570 75126 367606 77148
rect 527408 77140 527414 77148
rect 527466 77184 527472 77192
rect 527466 77148 527478 77184
rect 527466 77140 527472 77148
rect 526832 77100 526838 77108
rect 372190 77064 526838 77100
rect 372190 75112 372226 77064
rect 526832 77056 526838 77064
rect 526890 77100 526896 77108
rect 526890 77064 526898 77100
rect 526890 77056 526896 77064
rect 526472 77016 526478 77024
rect 376814 76980 526478 77016
rect 376814 75142 376850 76980
rect 526472 76972 526478 76980
rect 526530 76972 526536 77024
rect 525320 76932 525326 76942
rect 381442 76896 525326 76932
rect 381442 75134 381478 76896
rect 525320 76890 525326 76896
rect 525378 76932 525384 76942
rect 525378 76896 525386 76932
rect 525378 76890 525384 76896
rect 527192 76848 527198 76856
rect 390702 76812 527198 76848
rect 390702 75114 390738 76812
rect 527192 76804 527198 76812
rect 527250 76848 527256 76856
rect 527250 76812 527258 76848
rect 527250 76804 527256 76812
rect 527048 76764 527054 76772
rect 395330 76728 527054 76764
rect 395330 75126 395366 76728
rect 527048 76720 527054 76728
rect 527106 76764 527112 76772
rect 527106 76728 527114 76764
rect 527106 76720 527112 76728
rect 526688 76680 526694 76688
rect 399936 76644 526694 76680
rect 399936 75150 399972 76644
rect 526688 76636 526694 76644
rect 526746 76680 526752 76688
rect 526746 76644 526756 76680
rect 526746 76636 526752 76644
rect 525752 76596 525758 76604
rect 404574 76560 525758 76596
rect 404574 75172 404610 76560
rect 525752 76552 525758 76560
rect 525810 76596 525816 76604
rect 525810 76560 525820 76596
rect 525810 76552 525816 76560
rect 527336 76512 527342 76520
rect 413822 76476 527342 76512
rect 413822 75128 413858 76476
rect 527336 76468 527342 76476
rect 527394 76512 527400 76520
rect 527394 76476 527404 76512
rect 527394 76468 527400 76476
rect 526760 76428 526766 76436
rect 418462 76392 526766 76428
rect 418462 75136 418498 76392
rect 526760 76384 526766 76392
rect 526818 76384 526824 76436
rect 526400 76344 526406 76352
rect 423082 76308 526406 76344
rect 423082 75134 423118 76308
rect 526400 76300 526406 76308
rect 526458 76344 526464 76352
rect 526458 76308 526468 76344
rect 526458 76300 526464 76308
rect 525248 76260 525254 76268
rect 427710 76224 525254 76260
rect 427710 75168 427746 76224
rect 525248 76216 525254 76224
rect 525306 76260 525312 76268
rect 525306 76224 525314 76260
rect 525306 76216 525312 76224
rect 527120 76176 527126 76186
rect 436948 76140 527126 76176
rect 436948 75110 436984 76140
rect 527120 76134 527126 76140
rect 527178 76176 527184 76186
rect 527178 76140 527186 76176
rect 527178 76134 527184 76140
rect 526976 76092 526982 76100
rect 441602 76056 526982 76092
rect 441602 75138 441638 76056
rect 526976 76048 526982 76056
rect 527034 76092 527040 76100
rect 527034 76056 527042 76092
rect 527034 76048 527040 76056
rect 526616 76008 526622 76016
rect 446202 75972 526622 76008
rect 446202 75140 446238 75972
rect 526616 75964 526622 75972
rect 526674 76008 526680 76016
rect 526674 75972 526686 76008
rect 526674 75964 526680 75972
rect 525680 75924 525686 75934
rect 450838 75888 525686 75924
rect 450838 75146 450874 75888
rect 525680 75882 525686 75888
rect 525738 75924 525744 75934
rect 525738 75888 525748 75924
rect 525738 75882 525744 75888
rect 524816 75840 524822 75848
rect 460082 75804 524822 75840
rect 460082 75134 460118 75804
rect 524816 75796 524822 75804
rect 524874 75840 524880 75848
rect 524874 75804 524888 75840
rect 524874 75796 524880 75804
rect 525032 75756 525038 75764
rect 464706 75720 525038 75756
rect 464706 75156 464742 75720
rect 525032 75712 525038 75720
rect 525090 75756 525096 75764
rect 525090 75720 525098 75756
rect 525090 75712 525096 75720
rect 526328 75672 526334 75680
rect 469340 75636 526334 75672
rect 469340 75152 469376 75636
rect 526328 75628 526334 75636
rect 526386 75672 526392 75680
rect 526386 75636 526394 75672
rect 526386 75628 526392 75636
rect 525608 75588 525614 75596
rect 478598 75552 525614 75588
rect 478598 75138 478634 75552
rect 525608 75544 525614 75552
rect 525666 75588 525672 75596
rect 525666 75552 525680 75588
rect 525666 75544 525672 75552
rect 526904 75504 526910 75514
rect 483226 75468 526910 75504
rect 483226 75154 483262 75468
rect 526904 75462 526910 75468
rect 526962 75504 526968 75514
rect 526962 75468 526974 75504
rect 526962 75462 526968 75468
rect 525392 75420 525398 75428
rect 492462 75384 525398 75420
rect 492462 75126 492498 75384
rect 525392 75376 525398 75384
rect 525450 75420 525456 75428
rect 525450 75384 525460 75420
rect 525450 75376 525456 75384
rect 526544 75336 526550 75342
rect 497086 75300 526550 75336
rect 497088 75126 497124 75300
rect 526544 75290 526550 75300
rect 526602 75336 526608 75342
rect 526602 75300 526610 75336
rect 526602 75290 526608 75300
rect 215428 75100 215434 75109
rect 367549 69493 367831 69527
rect 367797 63382 367831 69493
rect 372172 69488 372472 69524
rect 376798 69492 377100 69528
rect 372436 63466 372472 69488
rect 377064 63550 377100 69492
rect 381430 69488 381726 69524
rect 381690 63634 381726 69488
rect 386054 69484 386346 69520
rect 390672 69488 390968 69524
rect 395300 69492 395612 69528
rect 386310 63718 386346 69484
rect 390932 63802 390968 69488
rect 395576 63886 395612 69492
rect 399928 69488 400218 69524
rect 404558 69488 404832 69524
rect 400182 63970 400218 69488
rect 404796 64054 404832 69488
rect 409180 69478 409466 69514
rect 413796 69492 414104 69528
rect 409430 64138 409466 69478
rect 414068 64222 414104 69492
rect 418426 69482 418730 69518
rect 418694 64306 418730 69482
rect 423066 69474 423356 69510
rect 427682 69488 427982 69524
rect 432312 69496 432602 69532
rect 436938 69496 437236 69532
rect 423320 64390 423356 69474
rect 427946 64474 427982 69488
rect 432566 64558 432602 69496
rect 437200 64642 437236 69496
rect 441548 69488 441866 69524
rect 446174 69496 446496 69532
rect 441830 64726 441866 69488
rect 446460 64810 446496 69496
rect 450818 69486 451114 69522
rect 455438 69500 455740 69536
rect 451078 64894 451114 69486
rect 455704 64978 455740 69500
rect 460064 69482 460370 69518
rect 464688 69486 465006 69522
rect 469310 69504 469624 69540
rect 460334 65062 460370 69482
rect 464970 65146 465006 69486
rect 469588 65230 469624 69504
rect 473944 69488 474248 69524
rect 478572 69498 478872 69534
rect 474212 65314 474248 69488
rect 478836 65398 478872 69498
rect 483200 69490 483502 69526
rect 487846 69490 488120 69526
rect 492428 69494 492752 69530
rect 497058 69502 497382 69538
rect 501694 69506 501990 69542
rect 483466 65482 483502 69490
rect 488084 65566 488120 69490
rect 492716 65650 492752 69494
rect 497346 65734 497382 69502
rect 501954 65818 501990 69506
rect 524168 65818 524174 65826
rect 501954 65782 524174 65818
rect 524168 65774 524174 65782
rect 524226 65818 524232 65826
rect 524226 65782 524236 65818
rect 524226 65774 524232 65782
rect 523664 65734 523670 65742
rect 497346 65698 523670 65734
rect 523664 65690 523670 65698
rect 523722 65734 523728 65742
rect 523722 65698 523736 65734
rect 523722 65690 523728 65698
rect 525824 65650 525830 65658
rect 492716 65614 525830 65650
rect 525824 65606 525830 65614
rect 525882 65650 525888 65658
rect 525882 65614 525896 65650
rect 525882 65606 525888 65614
rect 524456 65566 524462 65574
rect 488084 65530 524462 65566
rect 524456 65522 524462 65530
rect 524514 65566 524520 65574
rect 524514 65530 524530 65566
rect 524514 65522 524520 65530
rect 523952 65482 523958 65490
rect 483466 65446 523958 65482
rect 523952 65438 523958 65446
rect 524010 65482 524016 65490
rect 524010 65446 524022 65482
rect 524010 65438 524016 65446
rect 526112 65398 526118 65410
rect 478836 65362 526118 65398
rect 526112 65358 526118 65362
rect 526170 65398 526176 65410
rect 526170 65362 526184 65398
rect 526170 65358 526176 65362
rect 527264 65314 527270 65322
rect 474212 65278 527270 65314
rect 527264 65270 527270 65278
rect 527322 65314 527328 65322
rect 527322 65278 527336 65314
rect 527322 65270 527328 65278
rect 524240 65230 524246 65238
rect 469588 65194 524246 65230
rect 524240 65186 524246 65194
rect 524298 65230 524304 65238
rect 524298 65194 524310 65230
rect 524298 65186 524304 65194
rect 523736 65146 523742 65156
rect 464970 65110 523742 65146
rect 523736 65104 523742 65110
rect 523794 65146 523800 65156
rect 523794 65110 523806 65146
rect 523794 65104 523800 65110
rect 525896 65062 525902 65072
rect 460334 65026 525902 65062
rect 525896 65020 525902 65026
rect 525954 65062 525960 65072
rect 525954 65026 525966 65062
rect 525954 65020 525960 65026
rect 525464 64978 525470 64986
rect 455704 64942 525470 64978
rect 525464 64934 525470 64942
rect 525522 64978 525528 64986
rect 525522 64942 525534 64978
rect 525522 64934 525528 64942
rect 524672 64894 524678 64902
rect 451078 64858 524678 64894
rect 524672 64850 524678 64858
rect 524730 64894 524736 64902
rect 524730 64858 524740 64894
rect 524730 64850 524736 64858
rect 524528 64810 524534 64820
rect 446460 64774 524534 64810
rect 524528 64768 524534 64774
rect 524586 64810 524592 64820
rect 524586 64774 524600 64810
rect 524586 64768 524592 64774
rect 524024 64726 524030 64734
rect 441830 64690 524030 64726
rect 524024 64682 524030 64690
rect 524082 64726 524088 64734
rect 524082 64690 524094 64726
rect 524082 64682 524088 64690
rect 526184 64642 526190 64650
rect 437200 64606 526190 64642
rect 526184 64598 526190 64606
rect 526242 64642 526248 64650
rect 526242 64606 526252 64642
rect 526242 64598 526248 64606
rect 525104 64558 525110 64566
rect 432566 64522 525110 64558
rect 525104 64514 525110 64522
rect 525162 64558 525168 64566
rect 525162 64522 525176 64558
rect 525162 64514 525168 64522
rect 524888 64474 524894 64484
rect 427946 64438 524894 64474
rect 524888 64432 524894 64438
rect 524946 64474 524952 64484
rect 524946 64438 524958 64474
rect 524946 64432 524952 64438
rect 524312 64390 524318 64398
rect 423320 64354 524318 64390
rect 524312 64346 524318 64354
rect 524370 64390 524376 64398
rect 524370 64354 524380 64390
rect 524370 64346 524376 64354
rect 523808 64306 523814 64314
rect 418694 64270 523814 64306
rect 523808 64262 523814 64270
rect 523866 64306 523872 64314
rect 523866 64270 523882 64306
rect 523866 64262 523872 64270
rect 525968 64222 525974 64230
rect 414068 64186 525974 64222
rect 525968 64178 525974 64186
rect 526026 64222 526032 64230
rect 526026 64186 526038 64222
rect 526026 64178 526032 64186
rect 525536 64138 525542 64146
rect 409430 64102 525542 64138
rect 525536 64094 525542 64102
rect 525594 64138 525600 64146
rect 525594 64102 525604 64138
rect 525594 64094 525600 64102
rect 524744 64054 524750 64062
rect 404796 64018 524750 64054
rect 524744 64010 524750 64018
rect 524802 64054 524808 64062
rect 524802 64018 524816 64054
rect 524802 64010 524808 64018
rect 524600 63970 524606 63978
rect 400182 63934 524606 63970
rect 524600 63926 524606 63934
rect 524658 63970 524664 63978
rect 524658 63934 524668 63970
rect 524658 63926 524664 63934
rect 524096 63886 524102 63894
rect 395576 63850 524102 63886
rect 524096 63842 524102 63850
rect 524154 63886 524160 63894
rect 524154 63850 524166 63886
rect 524154 63842 524160 63850
rect 526256 63802 526262 63810
rect 390932 63766 526262 63802
rect 526256 63758 526262 63766
rect 526314 63802 526320 63810
rect 526314 63766 526324 63802
rect 526314 63758 526320 63766
rect 525176 63718 525182 63726
rect 386310 63682 525182 63718
rect 525176 63674 525182 63682
rect 525234 63718 525240 63726
rect 525234 63682 525248 63718
rect 525234 63674 525240 63682
rect 524960 63634 524966 63642
rect 381690 63598 524966 63634
rect 524960 63590 524966 63598
rect 525018 63634 525024 63642
rect 525018 63598 525030 63634
rect 525018 63590 525024 63598
rect 524384 63550 524390 63558
rect 377064 63514 524390 63550
rect 524384 63506 524390 63514
rect 524442 63550 524448 63558
rect 524442 63514 524454 63550
rect 524442 63506 524448 63514
rect 523880 63466 523886 63474
rect 372436 63430 523886 63466
rect 523880 63422 523886 63430
rect 523938 63466 523944 63474
rect 523938 63430 523946 63466
rect 523938 63422 523944 63430
rect 526040 63382 526046 63390
rect 367797 63348 526046 63382
rect 421972 63346 526046 63348
rect 526040 63338 526046 63346
rect 526098 63382 526104 63390
rect 526098 63346 526108 63382
rect 526098 63338 526104 63346
rect 385984 63241 385990 63293
rect 386042 63285 386048 63293
rect 544424 63285 544430 63292
rect 386042 63249 544430 63285
rect 386042 63241 386048 63249
rect 544424 63240 544430 63249
rect 544482 63285 544488 63292
rect 544482 63249 544497 63285
rect 544482 63240 544488 63249
rect 416036 63201 416042 63210
rect 416032 63165 416042 63201
rect 416036 63158 416042 63165
rect 416094 63201 416100 63210
rect 480545 63201 480551 63208
rect 416094 63165 480551 63201
rect 416094 63158 416100 63165
rect 480545 63156 480551 63165
rect 480603 63201 480609 63208
rect 544340 63201 544346 63208
rect 480603 63165 544346 63201
rect 480603 63156 480609 63165
rect 544340 63156 544346 63165
rect 544398 63201 544404 63208
rect 544398 63165 544413 63201
rect 544398 63156 544404 63165
rect 415952 63117 415958 63126
rect 415948 63081 415958 63117
rect 415952 63074 415958 63081
rect 416010 63117 416016 63126
rect 480629 63117 480635 63124
rect 416010 63081 480635 63117
rect 416010 63074 416016 63081
rect 480629 63072 480635 63081
rect 480687 63117 480693 63124
rect 544256 63117 544262 63124
rect 480687 63081 544262 63117
rect 480687 63072 480693 63081
rect 544256 63072 544262 63081
rect 544314 63117 544320 63124
rect 544314 63081 544329 63117
rect 544314 63072 544320 63081
rect 415868 63033 415874 63042
rect 415862 62997 415874 63033
rect 415868 62990 415874 62997
rect 415926 63033 415932 63042
rect 480713 63033 480719 63040
rect 415926 62997 480719 63033
rect 415926 62990 415932 62997
rect 480713 62988 480719 62997
rect 480771 63033 480777 63040
rect 544172 63033 544178 63040
rect 480771 62997 544178 63033
rect 480771 62988 480777 62997
rect 544172 62988 544178 62997
rect 544230 63033 544236 63040
rect 544230 62997 544245 63033
rect 544230 62988 544236 62997
rect 415784 62949 415790 62957
rect 415775 62913 415790 62949
rect 415784 62905 415790 62913
rect 415842 62949 415848 62957
rect 480797 62949 480803 62956
rect 415842 62913 480803 62949
rect 415842 62905 415848 62913
rect 480797 62904 480803 62913
rect 480855 62949 480861 62956
rect 544088 62949 544094 62956
rect 480855 62913 544094 62949
rect 480855 62904 480861 62913
rect 544088 62904 544094 62913
rect 544146 62949 544152 62956
rect 544146 62913 544161 62949
rect 544146 62904 544152 62913
rect 480881 62865 480887 62872
rect 480874 62829 480887 62865
rect 480881 62820 480887 62829
rect 480939 62865 480945 62872
rect 544004 62865 544010 62872
rect 480939 62829 544010 62865
rect 480939 62820 480945 62829
rect 544004 62820 544010 62829
rect 544062 62865 544068 62872
rect 544062 62829 544077 62865
rect 544062 62820 544068 62829
rect 480965 62781 480971 62788
rect 480958 62745 480971 62781
rect 480965 62736 480971 62745
rect 481023 62781 481029 62788
rect 543920 62781 543926 62788
rect 481023 62745 543926 62781
rect 481023 62736 481029 62745
rect 543920 62736 543926 62745
rect 543978 62781 543984 62788
rect 543978 62745 543993 62781
rect 543978 62736 543984 62745
rect 481049 62697 481055 62704
rect 481042 62661 481055 62697
rect 481049 62652 481055 62661
rect 481107 62697 481113 62704
rect 543836 62697 543842 62704
rect 481107 62661 543842 62697
rect 481107 62652 481113 62661
rect 543836 62652 543842 62661
rect 543894 62697 543900 62704
rect 543894 62661 543909 62697
rect 543894 62652 543900 62661
rect 481133 62613 481139 62620
rect 481126 62577 481139 62613
rect 481133 62568 481139 62577
rect 481191 62613 481197 62620
rect 543752 62613 543758 62620
rect 481191 62577 543758 62613
rect 481191 62568 481197 62577
rect 543752 62568 543758 62577
rect 543810 62613 543816 62620
rect 543810 62577 543825 62613
rect 543810 62568 543816 62577
rect 481217 62529 481223 62536
rect 481210 62493 481223 62529
rect 481217 62484 481223 62493
rect 481275 62529 481281 62536
rect 543668 62529 543674 62536
rect 481275 62493 543674 62529
rect 481275 62484 481281 62493
rect 543668 62484 543674 62493
rect 543726 62529 543732 62536
rect 543726 62493 543741 62529
rect 543726 62484 543732 62493
rect 481301 62445 481307 62452
rect 481294 62409 481307 62445
rect 481301 62400 481307 62409
rect 481359 62445 481365 62452
rect 543584 62445 543590 62452
rect 481359 62409 543590 62445
rect 481359 62400 481365 62409
rect 543584 62400 543590 62409
rect 543642 62445 543648 62452
rect 543642 62409 543657 62445
rect 543642 62400 543648 62409
rect 481385 62361 481391 62368
rect 481378 62325 481391 62361
rect 481385 62316 481391 62325
rect 481443 62361 481449 62368
rect 543500 62361 543506 62368
rect 481443 62325 543506 62361
rect 481443 62316 481449 62325
rect 543500 62316 543506 62325
rect 543558 62361 543564 62368
rect 543558 62325 543573 62361
rect 543558 62316 543564 62325
rect 481469 62277 481475 62284
rect 481462 62241 481475 62277
rect 481469 62232 481475 62241
rect 481527 62277 481533 62284
rect 543416 62277 543422 62284
rect 481527 62241 543422 62277
rect 481527 62232 481533 62241
rect 543416 62232 543422 62241
rect 543474 62277 543480 62284
rect 543474 62241 543489 62277
rect 543474 62232 543480 62241
rect 374007 62212 374013 62222
rect 373993 62176 374013 62212
rect 374007 62170 374013 62176
rect 374065 62212 374071 62222
rect 374065 62176 408736 62212
rect 481553 62193 481559 62200
rect 374065 62170 374071 62176
rect 374129 62128 374135 62138
rect 374112 62092 374135 62128
rect 374129 62086 374135 62092
rect 374187 62128 374193 62138
rect 374187 62092 408652 62128
rect 374187 62086 374193 62092
rect 291884 61975 408551 62049
rect 291884 61969 291958 61975
rect 83659 61744 83665 61969
rect 83739 61958 291958 61969
rect 83739 61906 84254 61958
rect 84306 61906 291958 61958
rect 83739 61895 291958 61906
rect 83739 61744 83745 61895
rect 292060 61889 292066 61941
rect 292118 61933 292124 61941
rect 292118 61897 408417 61933
rect 292118 61889 292124 61897
rect 292144 61805 292150 61857
rect 292202 61849 292208 61857
rect 292202 61813 408333 61849
rect 292202 61805 292208 61813
rect 340617 61765 340623 61774
rect 340615 61729 340623 61765
rect 340617 61722 340623 61729
rect 340675 61765 340681 61774
rect 340675 61729 408249 61765
rect 340675 61722 340681 61729
rect 340533 61681 340539 61690
rect 340528 61645 340539 61681
rect 340533 61638 340539 61645
rect 340591 61681 340597 61690
rect 340591 61645 408165 61681
rect 340591 61638 340597 61645
rect 240186 61565 290746 61601
rect 340449 61597 340455 61606
rect 240186 61371 240222 61565
rect 289935 61501 289941 61503
rect 282179 61465 289941 61501
rect 289935 61451 289941 61465
rect 289993 61451 289999 61503
rect 290019 61417 290025 61422
rect 282179 61381 290025 61417
rect 187227 61335 240222 61371
rect 290019 61370 290025 61381
rect 290077 61370 290083 61422
rect 183932 59797 185250 59846
rect 183932 59273 183998 59797
rect 185192 59273 185250 59797
rect 183932 59224 185250 59273
rect 83265 58763 83288 58815
rect 83340 58763 86020 58815
rect 185147 58346 186988 58427
rect 30168 57209 30174 57217
rect 30158 57173 30174 57209
rect 30168 57165 30174 57173
rect 30226 57209 30232 57217
rect 76398 57209 76404 57217
rect 30226 57173 76404 57209
rect 30226 57165 30232 57173
rect 76398 57165 76404 57173
rect 76456 57165 76462 57217
rect 29999 57125 30005 57133
rect 29991 57089 30005 57125
rect 29999 57081 30005 57089
rect 30057 57125 30063 57133
rect 70603 57125 70609 57133
rect 30057 57089 70609 57125
rect 30057 57081 30063 57089
rect 70603 57081 70609 57089
rect 70661 57081 70667 57133
rect 30083 57041 30089 57049
rect 30076 57005 30089 57041
rect 30083 56997 30089 57005
rect 30141 57041 30147 57049
rect 69962 57041 69968 57049
rect 30141 57005 69968 57041
rect 30141 56997 30147 57005
rect 69962 56997 69968 57005
rect 70020 56997 70026 57049
rect 31007 56957 31013 56965
rect 31003 56921 31013 56957
rect 31007 56913 31013 56921
rect 31065 56957 31071 56965
rect 67372 56957 67378 56965
rect 31065 56921 67378 56957
rect 31065 56913 31071 56921
rect 67372 56913 67378 56921
rect 67430 56913 67436 56965
rect 30840 56873 30846 56881
rect 30830 56837 30846 56873
rect 30840 56829 30846 56837
rect 30898 56873 30904 56881
rect 64927 56873 64933 56881
rect 30898 56837 64933 56873
rect 30898 56829 30904 56837
rect 64927 56829 64933 56837
rect 64985 56829 64991 56881
rect 9246 55843 9252 55895
rect 9304 55883 9310 55895
rect 9304 55855 12968 55883
rect 9304 55843 9310 55855
rect 9358 55716 9364 55768
rect 9416 55756 9422 55768
rect 9416 55728 12981 55756
rect 9416 55716 9422 55728
rect 9470 55611 9476 55663
rect 9528 55651 9534 55663
rect 9528 55623 12968 55651
rect 9528 55611 9534 55623
rect 9583 55536 9589 55545
rect 9582 55501 9589 55536
rect 9583 55493 9589 55501
rect 9641 55536 9647 55545
rect 9641 55501 12951 55536
rect 9641 55493 9647 55501
rect 184763 54407 186122 54490
rect 187227 54044 187263 61335
rect 289767 61333 289773 61341
rect 282178 61297 289773 61333
rect 289767 61289 289773 61297
rect 289825 61289 289831 61341
rect 289854 61249 289860 61257
rect 282176 61213 289860 61249
rect 289854 61205 289860 61213
rect 289912 61205 289918 61257
rect 290710 60908 290746 61565
rect 340444 61561 340455 61597
rect 340449 61554 340455 61561
rect 340507 61597 340513 61606
rect 340507 61561 408081 61597
rect 340507 61554 340513 61561
rect 292314 61471 292320 61523
rect 292372 61513 292378 61523
rect 292372 61477 407997 61513
rect 292372 61471 292378 61477
rect 292398 61385 292404 61437
rect 292456 61429 292462 61437
rect 292456 61393 407913 61429
rect 292456 61385 292462 61393
rect 292479 61301 292485 61353
rect 292537 61345 292543 61353
rect 292537 61309 407829 61345
rect 292537 61301 292543 61309
rect 292230 61218 292236 61270
rect 292288 61261 292294 61270
rect 292288 61225 407745 61261
rect 292288 61218 292294 61225
rect 374248 61133 374254 61185
rect 374306 61177 374312 61185
rect 374306 61141 407661 61177
rect 374306 61133 374312 61141
rect 341052 61093 341058 61125
rect 341049 61057 341058 61093
rect 341052 61025 341058 61057
rect 341158 61093 341164 61125
rect 341158 61057 407577 61093
rect 341158 61025 341164 61057
rect 391300 60956 391306 61008
rect 391358 61000 391364 61008
rect 391358 60964 407128 61000
rect 391358 60956 391364 60964
rect 290710 60872 407031 60908
rect 405582 59336 405782 60595
rect 405882 59336 406082 60595
rect 406182 59336 406382 60595
rect 406995 60170 407031 60872
rect 407092 60254 407128 60964
rect 407541 60422 407577 61057
rect 407625 60506 407661 61141
rect 407709 60674 407745 61225
rect 407793 60758 407829 61309
rect 407877 60842 407913 61393
rect 407961 60926 407997 61477
rect 408045 61010 408081 61561
rect 408129 61094 408165 61645
rect 408213 61178 408249 61729
rect 408297 61262 408333 61813
rect 408381 61346 408417 61897
rect 408477 61592 408551 61975
rect 408616 61689 408652 62092
rect 408700 61773 408736 62176
rect 481546 62157 481559 62193
rect 481553 62148 481559 62157
rect 481611 62193 481617 62200
rect 543332 62193 543338 62200
rect 481611 62157 543338 62193
rect 481611 62148 481617 62157
rect 543332 62148 543338 62157
rect 543390 62193 543396 62200
rect 543390 62157 543405 62193
rect 543390 62148 543396 62157
rect 481637 62109 481643 62116
rect 481630 62073 481643 62109
rect 481637 62064 481643 62073
rect 481695 62109 481701 62116
rect 543248 62109 543254 62116
rect 481695 62073 543254 62109
rect 481695 62064 481701 62073
rect 543248 62064 543254 62073
rect 543306 62109 543312 62116
rect 543306 62073 543321 62109
rect 543306 62064 543312 62073
rect 481721 62025 481727 62032
rect 481714 61989 481727 62025
rect 481721 61980 481727 61989
rect 481779 62025 481785 62032
rect 543164 62025 543170 62032
rect 481779 61989 543170 62025
rect 481779 61980 481785 61989
rect 543164 61980 543170 61989
rect 543222 62025 543228 62032
rect 543222 61989 543237 62025
rect 543222 61980 543228 61989
rect 481805 61941 481811 61948
rect 481798 61905 481811 61941
rect 481805 61896 481811 61905
rect 481863 61941 481869 61948
rect 543080 61941 543086 61948
rect 481863 61905 543086 61941
rect 481863 61896 481869 61905
rect 543080 61896 543086 61905
rect 543138 61941 543144 61948
rect 543138 61905 543153 61941
rect 543138 61896 543144 61905
rect 415700 61857 415706 61864
rect 415695 61821 415706 61857
rect 415700 61812 415706 61821
rect 415758 61857 415764 61864
rect 542996 61857 543002 61864
rect 415758 61821 543002 61857
rect 415758 61812 415764 61821
rect 542996 61812 543002 61821
rect 543054 61857 543060 61864
rect 543054 61821 543069 61857
rect 543054 61812 543060 61821
rect 542912 61773 542918 61780
rect 408700 61737 542918 61773
rect 542912 61728 542918 61737
rect 542970 61773 542976 61780
rect 542970 61737 542985 61773
rect 542970 61728 542976 61737
rect 542828 61689 542834 61696
rect 408616 61653 542834 61689
rect 542828 61644 542834 61653
rect 542886 61689 542892 61696
rect 542886 61653 542901 61689
rect 542886 61644 542892 61653
rect 432532 61624 522382 61625
rect 430744 61622 522382 61624
rect 408477 61588 430208 61592
rect 408477 61522 429774 61588
rect 430184 61522 430208 61588
rect 430744 61564 430758 61622
rect 431270 61607 522382 61622
rect 431270 61564 522319 61607
rect 430744 61560 522319 61564
rect 408477 61518 430208 61522
rect 430711 61514 430717 61522
rect 430706 61478 430717 61514
rect 430711 61470 430717 61478
rect 430769 61514 430775 61522
rect 522209 61514 522215 61523
rect 430769 61478 522215 61514
rect 430769 61470 430775 61478
rect 522209 61471 522215 61478
rect 522267 61514 522273 61523
rect 522267 61478 522277 61514
rect 522267 61471 522273 61478
rect 430794 61430 430800 61438
rect 430793 61394 430800 61430
rect 430794 61386 430800 61394
rect 430852 61430 430858 61438
rect 522125 61430 522131 61438
rect 430852 61394 522131 61430
rect 430852 61386 430858 61394
rect 522125 61386 522131 61394
rect 522183 61430 522189 61438
rect 522183 61394 522192 61430
rect 522306 61400 522319 61560
rect 522313 61395 522319 61400
rect 522371 61400 522382 61607
rect 522371 61395 522377 61400
rect 522183 61386 522189 61394
rect 542744 61346 542750 61354
rect 408381 61310 542750 61346
rect 542744 61302 542750 61310
rect 542802 61302 542808 61354
rect 565930 61289 567363 61773
rect 542660 61262 542666 61270
rect 408297 61226 542666 61262
rect 542660 61218 542666 61226
rect 542718 61262 542724 61270
rect 542718 61226 542733 61262
rect 542718 61218 542724 61226
rect 542576 61178 542582 61186
rect 408213 61142 542582 61178
rect 542576 61134 542582 61142
rect 542634 61178 542640 61186
rect 542634 61142 542649 61178
rect 542634 61134 542640 61142
rect 542492 61094 542498 61102
rect 408129 61058 542498 61094
rect 542492 61050 542498 61058
rect 542550 61094 542556 61102
rect 542550 61058 542565 61094
rect 542550 61050 542556 61058
rect 485622 61010 485628 61018
rect 408045 60974 485628 61010
rect 485622 60966 485628 60974
rect 485680 60966 485686 61018
rect 519074 61010 519080 61018
rect 519072 60974 519080 61010
rect 519074 60966 519080 60974
rect 519132 61010 519138 61018
rect 542408 61010 542414 61018
rect 519132 60974 542414 61010
rect 519132 60966 519138 60974
rect 542408 60966 542414 60974
rect 542466 61010 542472 61018
rect 542466 60974 542481 61010
rect 542466 60966 542472 60974
rect 485706 60926 485712 60934
rect 407961 60890 485712 60926
rect 485706 60882 485712 60890
rect 485764 60882 485770 60934
rect 518990 60882 518996 60934
rect 519048 60926 519054 60934
rect 542324 60926 542330 60934
rect 519048 60890 542330 60926
rect 519048 60882 519054 60890
rect 542324 60882 542330 60890
rect 542382 60926 542388 60934
rect 542382 60890 542397 60926
rect 542382 60882 542388 60890
rect 485788 60842 485794 60850
rect 407877 60806 485794 60842
rect 485788 60798 485794 60806
rect 485846 60798 485852 60850
rect 518906 60842 518912 60850
rect 518902 60806 518912 60842
rect 518906 60798 518912 60806
rect 518964 60842 518970 60850
rect 542240 60842 542246 60850
rect 518964 60806 542246 60842
rect 518964 60798 518970 60806
rect 542240 60798 542246 60806
rect 542298 60842 542304 60850
rect 542298 60806 542313 60842
rect 542298 60798 542304 60806
rect 485876 60758 485882 60766
rect 407793 60722 485882 60758
rect 485876 60714 485882 60722
rect 485934 60714 485940 60766
rect 518822 60758 518828 60766
rect 518816 60722 518828 60758
rect 518822 60714 518828 60722
rect 518880 60758 518886 60766
rect 542156 60758 542162 60766
rect 518880 60722 542162 60758
rect 518880 60714 518886 60722
rect 542156 60714 542162 60722
rect 542214 60758 542220 60766
rect 542214 60722 542229 60758
rect 542214 60714 542220 60722
rect 562701 60715 564300 61071
rect 485962 60674 485968 60682
rect 407709 60638 485968 60674
rect 485962 60630 485968 60638
rect 486020 60630 486026 60682
rect 518738 60674 518744 60682
rect 518730 60638 518744 60674
rect 518738 60630 518744 60638
rect 518796 60674 518802 60682
rect 542072 60674 542078 60682
rect 518796 60638 542078 60674
rect 518796 60630 518802 60638
rect 542072 60630 542078 60638
rect 542130 60674 542136 60682
rect 542130 60638 542145 60674
rect 562697 60665 564300 60715
rect 542130 60630 542136 60638
rect 481931 60590 481937 60599
rect 481923 60554 481937 60590
rect 481931 60547 481937 60554
rect 481989 60590 481995 60599
rect 486040 60590 486046 60598
rect 481989 60554 486046 60590
rect 481989 60547 481995 60554
rect 486040 60546 486046 60554
rect 486098 60546 486104 60598
rect 518654 60590 518660 60598
rect 518650 60554 518660 60590
rect 518654 60546 518660 60554
rect 518712 60590 518718 60598
rect 541988 60590 541994 60598
rect 518712 60554 541994 60590
rect 518712 60546 518718 60554
rect 541988 60546 541994 60554
rect 542046 60590 542052 60598
rect 542046 60554 542061 60590
rect 542046 60546 542052 60554
rect 486130 60506 486136 60514
rect 407625 60470 486136 60506
rect 486130 60462 486136 60470
rect 486188 60462 486194 60514
rect 518570 60506 518576 60514
rect 518566 60470 518576 60506
rect 518570 60462 518576 60470
rect 518628 60506 518634 60514
rect 541904 60506 541910 60514
rect 518628 60470 541910 60506
rect 518628 60462 518634 60470
rect 541904 60462 541910 60470
rect 541962 60506 541968 60514
rect 541962 60470 541977 60506
rect 561004 60504 561010 60512
rect 541962 60462 541968 60470
rect 557343 60458 558215 60494
rect 560987 60468 561010 60504
rect 561004 60460 561010 60468
rect 561062 60504 561068 60512
rect 561062 60468 561912 60504
rect 561062 60460 561068 60468
rect 486210 60422 486216 60430
rect 407541 60386 486216 60422
rect 486210 60378 486216 60386
rect 486268 60378 486274 60430
rect 518486 60422 518492 60430
rect 518478 60386 518492 60422
rect 518486 60378 518492 60386
rect 518544 60422 518550 60430
rect 541820 60422 541826 60430
rect 518544 60386 541826 60422
rect 518544 60378 518550 60386
rect 541820 60378 541826 60386
rect 541878 60422 541884 60430
rect 541878 60386 541893 60422
rect 541878 60378 541884 60386
rect 544416 60378 547288 60418
rect 422507 60338 422513 60346
rect 422493 60302 422513 60338
rect 422507 60294 422513 60302
rect 422565 60338 422571 60346
rect 486292 60338 486298 60346
rect 422565 60302 486298 60338
rect 422565 60294 422571 60302
rect 486292 60294 486298 60302
rect 486350 60294 486356 60346
rect 518402 60338 518408 60346
rect 518398 60302 518408 60338
rect 518402 60294 518408 60302
rect 518460 60338 518466 60346
rect 541736 60338 541742 60346
rect 518460 60302 541742 60338
rect 518460 60294 518466 60302
rect 541736 60294 541742 60302
rect 541794 60338 541800 60346
rect 541794 60302 541809 60338
rect 541794 60294 541800 60302
rect 486376 60254 486382 60262
rect 407092 60218 486382 60254
rect 486376 60210 486382 60218
rect 486434 60210 486440 60262
rect 518318 60254 518324 60262
rect 518312 60218 518324 60254
rect 518318 60210 518324 60218
rect 518376 60254 518382 60262
rect 541652 60254 541658 60262
rect 518376 60218 541658 60254
rect 518376 60210 518382 60218
rect 541652 60210 541658 60218
rect 541710 60254 541716 60262
rect 541710 60218 541725 60254
rect 541710 60210 541716 60218
rect 406995 60169 485594 60170
rect 486462 60169 486468 60178
rect 406995 60135 486468 60169
rect 406995 60134 485594 60135
rect 486462 60126 486468 60135
rect 486520 60126 486526 60178
rect 518234 60170 518240 60178
rect 518226 60134 518240 60170
rect 518234 60126 518240 60134
rect 518292 60170 518298 60178
rect 541568 60170 541574 60178
rect 518292 60134 541574 60170
rect 518292 60126 518298 60134
rect 541568 60126 541574 60134
rect 541626 60170 541632 60178
rect 541626 60134 541641 60170
rect 541626 60126 541632 60134
rect 406677 59916 407807 59944
rect 406677 59791 406725 59916
rect 406482 59616 406725 59791
rect 407761 59616 407807 59916
rect 406482 59583 407807 59616
rect 342744 58606 342790 59266
rect 342918 58606 343302 59266
rect 343430 58606 343814 59266
rect 343942 58606 344326 59266
rect 344454 58606 344838 59266
rect 344966 58606 345350 59266
rect 345478 58606 345862 59266
rect 345990 58606 346374 59266
rect 346502 58606 346886 59266
rect 347014 58606 347398 59266
rect 347526 58606 348422 59266
rect 348550 58606 348934 59266
rect 349062 58606 349446 59266
rect 349574 58606 349958 59266
rect 350086 58606 350470 59266
rect 350598 58606 350982 59266
rect 351110 58606 351494 59266
rect 351622 59265 353480 59266
rect 351622 59225 354006 59265
rect 351622 58638 352180 59225
rect 353960 58638 354006 59225
rect 406482 59165 406682 59583
rect 364620 58778 372098 58896
rect 351622 58606 354006 58638
rect 352133 58603 354006 58606
rect 364068 58418 370476 58536
rect 370358 57999 370476 58418
rect 371980 58014 372098 58778
rect 288004 56803 288010 56811
rect 282223 56767 288010 56803
rect 288004 56759 288010 56767
rect 288062 56759 288068 56811
rect 288504 56719 288510 56727
rect 282219 56683 288510 56719
rect 288504 56675 288510 56683
rect 288562 56675 288568 56727
rect 289182 56635 289188 56643
rect 282221 56599 289188 56635
rect 289182 56591 289188 56599
rect 289240 56591 289246 56643
rect 354356 54468 354362 54476
rect 351516 54432 354362 54468
rect 354356 54424 354362 54432
rect 354414 54424 354420 54476
rect 354370 54370 354406 54424
rect 186235 54012 186242 54020
rect 184738 53976 186242 54012
rect 186235 53968 186242 53976
rect 186294 53968 186301 54020
rect 187227 54008 187461 54044
rect 187135 53487 187495 53595
rect 184818 53382 186923 53465
rect 187135 52978 187243 53487
rect 184777 52870 187243 52978
rect 83362 52496 83370 52548
rect 83422 52496 86018 52548
rect 182377 52464 184035 52741
rect 184777 52549 184885 52870
rect 186469 52604 187820 52655
rect 186469 52451 186566 52604
rect 186479 52384 186566 52451
rect 187774 52384 187820 52604
rect 186479 52333 187820 52384
rect 287830 52170 287836 52178
rect 249595 52115 249601 52167
rect 249653 52155 249659 52167
rect 249653 52119 254703 52155
rect 282218 52134 287836 52170
rect 287830 52126 287836 52134
rect 287888 52126 287894 52178
rect 249653 52115 249659 52119
rect 288678 52086 288684 52094
rect 282207 52050 288684 52086
rect 288678 52042 288684 52050
rect 288736 52042 288742 52094
rect 248167 51956 248173 52008
rect 248225 51997 248231 52008
rect 289350 52002 289356 52010
rect 248225 51961 254734 51997
rect 282212 51966 289356 52002
rect 248225 51956 248231 51961
rect 289350 51958 289356 51966
rect 289408 51958 289414 52010
rect 248671 51866 248677 51918
rect 248729 51913 248735 51918
rect 248729 51877 254715 51913
rect 248729 51866 248735 51877
rect 249427 51786 249433 51838
rect 249485 51829 249491 51838
rect 249485 51793 254695 51829
rect 249485 51786 249491 51793
rect 248923 51661 248929 51713
rect 248981 51705 248987 51713
rect 250541 51705 250547 51717
rect 248981 51669 250547 51705
rect 248981 51661 248987 51669
rect 250541 51665 250547 51669
rect 250599 51665 250605 51717
rect 241588 51575 241594 51627
rect 241646 51619 241652 51627
rect 249763 51619 249769 51627
rect 241646 51583 249769 51619
rect 241646 51575 241652 51583
rect 249763 51575 249769 51583
rect 249821 51575 249827 51627
rect 241889 51432 241895 51484
rect 241947 51480 241953 51484
rect 249847 51480 249853 51488
rect 241947 51444 249853 51480
rect 241947 51432 241953 51444
rect 249847 51436 249853 51444
rect 249905 51436 249911 51488
rect 241504 51305 241510 51357
rect 241562 51345 241568 51357
rect 249931 51345 249937 51354
rect 241562 51317 249937 51345
rect 241562 51305 241568 51317
rect 249931 51302 249937 51317
rect 249989 51302 249995 51354
rect 246013 51140 246019 51192
rect 246071 51184 246077 51192
rect 248001 51184 248007 51192
rect 246071 51148 248007 51184
rect 246071 51140 246077 51148
rect 248001 51140 248007 51148
rect 248059 51140 248065 51192
rect 241176 51074 241228 51080
rect 250016 51062 250022 51074
rect 241228 51034 250022 51062
rect 250016 51022 250022 51034
rect 250074 51022 250080 51074
rect 241176 51016 241228 51022
rect 9022 49934 9028 49986
rect 9080 49974 9086 49986
rect 9080 49946 12957 49974
rect 9080 49934 9086 49946
rect 522293 49906 522299 50114
rect 9134 49824 9140 49876
rect 9192 49864 9198 49876
rect 522289 49870 522299 49906
rect 9192 49836 12987 49864
rect 522293 49862 522299 49870
rect 522351 49930 522357 50114
rect 530286 50048 530326 50642
rect 530398 50188 530438 50658
rect 536186 50334 536226 50642
rect 536326 50462 536366 50636
rect 536326 50422 541828 50462
rect 536186 50294 541708 50334
rect 530398 50148 541588 50188
rect 530286 50008 541468 50048
rect 540268 49930 540337 49931
rect 522351 49920 540337 49930
rect 522351 49870 540273 49920
rect 522351 49862 522357 49870
rect 354278 49836 354284 49844
rect 9192 49824 9198 49836
rect 351476 49800 354284 49836
rect 354278 49792 354284 49800
rect 354336 49792 354342 49844
rect 522209 49822 522215 49830
rect 522205 49786 522215 49822
rect 522209 49778 522215 49786
rect 522267 49822 522273 49830
rect 540158 49822 540164 49836
rect 522267 49786 540164 49822
rect 522267 49778 522273 49786
rect 540158 49784 540164 49786
rect 540216 49784 540222 49836
rect 8798 49697 8804 49749
rect 8856 49737 8862 49749
rect 522125 49738 522131 49745
rect 8856 49709 13003 49737
rect 8856 49697 8862 49709
rect 522121 49702 522131 49738
rect 522125 49693 522131 49702
rect 522183 49738 522189 49745
rect 540046 49738 540052 49751
rect 522183 49702 540052 49738
rect 522183 49693 522189 49702
rect 540046 49699 540052 49702
rect 540104 49699 540110 49751
rect 540268 49693 540273 49870
rect 540332 49693 540337 49920
rect 540268 49687 540337 49693
rect 8910 49581 8916 49633
rect 8968 49621 8974 49633
rect 8968 49593 12967 49621
rect 8968 49581 8974 49593
rect 365279 48708 365359 49138
rect 371987 48812 372023 49330
rect 372930 48917 372966 49307
rect 374007 48917 374013 48925
rect 372930 48881 374013 48917
rect 374007 48873 374013 48881
rect 374065 48873 374071 48925
rect 374129 48812 374135 48820
rect 371987 48776 374135 48812
rect 374129 48768 374135 48776
rect 374187 48768 374193 48820
rect 374248 48708 374254 48716
rect 365279 48672 374254 48708
rect 374248 48664 374254 48672
rect 374306 48664 374312 48716
rect 422508 47562 422514 47570
rect 248076 47493 248082 47545
rect 248134 47537 248140 47545
rect 287923 47537 287929 47545
rect 248134 47501 254908 47537
rect 282219 47501 287929 47537
rect 248134 47493 248140 47501
rect 287923 47493 287929 47501
rect 287981 47493 287987 47545
rect 420993 47526 422514 47562
rect 422508 47518 422514 47526
rect 422566 47518 422572 47570
rect 249003 47409 249009 47461
rect 249061 47453 249067 47461
rect 288422 47453 288428 47461
rect 249061 47417 254902 47453
rect 282218 47417 288428 47453
rect 249061 47409 249067 47417
rect 288422 47409 288428 47417
rect 288480 47409 288486 47461
rect 249681 47325 249687 47377
rect 249739 47369 249745 47377
rect 289097 47369 289103 47377
rect 249739 47333 254893 47369
rect 282207 47333 289103 47369
rect 249739 47325 249745 47333
rect 289097 47325 289103 47333
rect 289155 47325 289161 47377
rect 541428 47342 541468 50008
rect 541548 47462 541588 50148
rect 541668 47582 541708 50294
rect 541788 47702 541828 50422
rect 544416 47862 544456 60378
rect 557254 60346 558101 60382
rect 544496 60258 547364 60298
rect 544496 47942 544536 60258
rect 557202 60234 558012 60270
rect 544576 60138 547436 60178
rect 544576 48022 544616 60138
rect 557127 60122 557924 60158
rect 544656 60018 547512 60058
rect 552682 60042 555620 60078
rect 544656 48102 544696 60018
rect 552608 59930 555530 59966
rect 552536 59838 555444 59874
rect 552470 59746 555230 59782
rect 555194 59622 555230 59746
rect 555408 59694 555444 59838
rect 555494 59766 555530 59930
rect 555584 59838 555620 60042
rect 557888 59910 557924 60122
rect 557976 59982 558012 60234
rect 558065 60054 558101 60346
rect 558179 60126 558215 60458
rect 562697 60236 562759 60665
rect 564261 60236 564300 60665
rect 561920 60220 561926 60228
rect 561578 60184 561926 60220
rect 561920 60176 561926 60184
rect 561978 60220 561984 60228
rect 561978 60184 561990 60220
rect 561978 60176 561984 60184
rect 562697 60167 564300 60236
rect 562402 60138 562408 60146
rect 561244 60126 561250 60134
rect 558179 60090 561250 60126
rect 561244 60082 561250 60090
rect 561302 60126 561308 60134
rect 561302 60090 561310 60126
rect 561572 60102 562408 60138
rect 562402 60094 562408 60102
rect 562460 60138 562466 60146
rect 562460 60102 562478 60138
rect 562460 60094 562466 60102
rect 561302 60082 561308 60090
rect 562042 60054 562048 60062
rect 558065 60018 562048 60054
rect 562042 60010 562048 60018
rect 562100 60054 562106 60062
rect 562100 60018 562118 60054
rect 562100 60010 562106 60018
rect 562640 59982 562646 59990
rect 557976 59946 562646 59982
rect 562640 59938 562646 59946
rect 562698 59938 562704 59990
rect 564795 59910 564801 59918
rect 557888 59874 564801 59910
rect 564795 59866 564801 59874
rect 564853 59866 564859 59918
rect 561122 59838 561128 59846
rect 555584 59802 561128 59838
rect 561122 59794 561128 59802
rect 561180 59838 561186 59846
rect 561180 59802 561194 59838
rect 561180 59794 561186 59802
rect 561684 59766 561690 59774
rect 555494 59730 561690 59766
rect 561684 59722 561690 59730
rect 561742 59766 561748 59774
rect 561742 59730 561754 59766
rect 561742 59722 561748 59730
rect 562162 59694 562168 59702
rect 555408 59658 562168 59694
rect 562162 59650 562168 59658
rect 562220 59694 562226 59702
rect 562220 59658 562232 59694
rect 562220 59650 562226 59658
rect 562522 59622 562528 59630
rect 555194 59586 562528 59622
rect 562522 59578 562528 59586
rect 562580 59622 562586 59630
rect 562580 59586 562594 59622
rect 562580 59578 562586 59586
rect 566879 58998 567363 61289
rect 565173 58968 567363 58998
rect 565173 58543 565210 58968
rect 566611 58543 567363 58968
rect 565173 58514 567363 58543
rect 562996 58210 567778 58250
rect 563118 58090 567900 58130
rect 563232 57970 568016 58010
rect 563338 57850 568138 57890
rect 563458 57730 568264 57770
rect 563574 57610 568374 57650
rect 563680 57490 568496 57530
rect 563790 57370 568614 57410
rect 563908 57250 568736 57290
rect 564018 57130 568858 57170
rect 564128 57010 568982 57050
rect 564238 56890 569106 56930
rect 564354 56770 569222 56810
rect 564458 56650 569344 56690
rect 564570 56530 569458 56570
rect 564680 56410 569572 56450
rect 568602 54658 568608 54670
rect 560792 54630 568608 54658
rect 568602 54618 568608 54630
rect 568660 54618 568666 54670
rect 568718 54538 568724 54550
rect 560766 54510 568724 54538
rect 568718 54498 568724 54510
rect 568776 54498 568782 54550
rect 567706 54408 567712 54420
rect 560750 54380 567712 54408
rect 567706 54368 567712 54380
rect 567764 54368 567770 54420
rect 567818 54300 567824 54312
rect 560766 54272 567824 54300
rect 567818 54260 567824 54272
rect 567876 54260 567882 54312
rect 567482 48750 567488 48762
rect 560758 48722 567488 48750
rect 567482 48710 567488 48722
rect 567540 48710 567546 48762
rect 567594 48636 567600 48648
rect 560788 48608 567600 48636
rect 567594 48596 567600 48608
rect 567652 48596 567658 48648
rect 567258 48510 567264 48522
rect 560716 48482 567264 48510
rect 567258 48470 567264 48482
rect 567316 48470 567322 48522
rect 567370 48386 567376 48398
rect 560774 48358 567376 48386
rect 567370 48346 567376 48358
rect 567428 48346 567434 48398
rect 561564 48102 561570 48108
rect 544656 48062 561570 48102
rect 561564 48056 561570 48062
rect 561622 48056 561628 48108
rect 562282 48022 562288 48028
rect 544576 47982 562288 48022
rect 562282 47976 562288 47982
rect 562340 47976 562346 48028
rect 562764 47942 562770 47948
rect 544496 47902 562770 47942
rect 562764 47896 562770 47902
rect 562822 47896 562828 47948
rect 562880 47862 562886 47868
rect 544416 47822 562886 47862
rect 562880 47816 562886 47822
rect 562938 47816 562944 47868
rect 560956 47702 560962 47708
rect 541788 47662 560962 47702
rect 560956 47656 560962 47662
rect 561014 47656 561020 47708
rect 561082 47582 561088 47594
rect 541668 47542 561088 47582
rect 561140 47542 561146 47594
rect 560716 47462 560722 47468
rect 541548 47422 560722 47462
rect 560716 47416 560722 47422
rect 560774 47416 560780 47468
rect 560838 47342 560844 47348
rect 541428 47302 560844 47342
rect 560838 47296 560844 47302
rect 560896 47296 560902 47348
rect 420754 47158 421778 47190
rect 541584 47176 567994 47184
rect 420754 47148 421781 47158
rect 420754 47023 420803 47148
rect 421743 47023 421781 47148
rect 420754 46988 421781 47023
rect 541584 47124 567936 47176
rect 567988 47124 567994 47176
rect 83454 46896 83460 46897
rect 83452 46846 83460 46896
rect 83454 46845 83460 46846
rect 83512 46896 83518 46897
rect 83512 46846 86047 46896
rect 83512 46845 83518 46846
rect 403880 46464 404079 46486
rect 402560 45630 402760 46056
rect 403120 45712 403156 46089
rect 403386 45797 403422 46162
rect 403663 45888 403699 46188
rect 403880 46006 403905 46464
rect 404057 46006 404079 46464
rect 403880 45980 404079 46006
rect 404186 46458 404385 46486
rect 404186 46000 404206 46458
rect 404358 46000 404385 46458
rect 420747 46173 421736 46211
rect 420747 46034 420789 46173
rect 421670 46034 421736 46173
rect 420747 46003 421736 46034
rect 404186 45980 404385 46000
rect 415700 45888 415706 45896
rect 403663 45852 415706 45888
rect 415700 45844 415706 45852
rect 415758 45888 415764 45896
rect 415758 45852 415771 45888
rect 415758 45844 415764 45852
rect 415784 45797 415790 45805
rect 403386 45761 415790 45797
rect 415784 45753 415790 45761
rect 415842 45797 415848 45805
rect 415842 45761 415857 45797
rect 415842 45753 415848 45761
rect 415868 45712 415874 45719
rect 403120 45676 415874 45712
rect 415868 45667 415874 45676
rect 415926 45712 415932 45719
rect 415926 45676 415937 45712
rect 415926 45667 415932 45676
rect 353766 45204 353772 45212
rect 351490 45168 353772 45204
rect 353766 45160 353772 45168
rect 353824 45160 353830 45212
rect 391650 45018 391672 45630
rect 392309 45018 402760 45630
rect 402906 45622 402958 45628
rect 415952 45614 415958 45621
rect 402958 45578 415958 45614
rect 402906 45564 402958 45570
rect 415952 45569 415958 45578
rect 416010 45614 416016 45621
rect 416010 45578 416018 45614
rect 416010 45569 416016 45578
rect 402908 45515 402960 45521
rect 416036 45508 416042 45514
rect 402960 45472 416042 45508
rect 402908 45457 402960 45463
rect 416036 45462 416042 45472
rect 416094 45508 416100 45514
rect 416094 45472 416102 45508
rect 416094 45462 416100 45472
rect 452721 44756 452727 44764
rect 452712 44720 452727 44756
rect 452721 44712 452727 44720
rect 452779 44756 452785 44764
rect 480545 44756 480551 44761
rect 452779 44720 480551 44756
rect 452779 44712 452785 44720
rect 480545 44709 480551 44720
rect 480603 44756 480609 44761
rect 480603 44720 480617 44756
rect 480603 44709 480609 44720
rect 446714 44672 446720 44680
rect 446698 44636 446720 44672
rect 446714 44628 446720 44636
rect 446772 44672 446778 44680
rect 480629 44672 480635 44677
rect 446772 44636 480635 44672
rect 446772 44628 446778 44636
rect 480629 44625 480635 44636
rect 480687 44672 480693 44677
rect 480687 44636 480701 44672
rect 480687 44625 480693 44636
rect 452559 44588 452565 44596
rect 452550 44552 452565 44588
rect 452559 44544 452565 44552
rect 452617 44588 452623 44596
rect 480713 44588 480719 44593
rect 452617 44552 480719 44588
rect 452617 44544 452623 44552
rect 480713 44541 480719 44552
rect 480771 44588 480777 44593
rect 480771 44552 480785 44588
rect 480771 44541 480777 44552
rect 446878 44504 446884 44512
rect 446862 44468 446884 44504
rect 446878 44460 446884 44468
rect 446936 44504 446942 44512
rect 480797 44504 480803 44509
rect 446936 44468 480803 44504
rect 446936 44460 446942 44468
rect 480797 44457 480803 44468
rect 480855 44504 480861 44509
rect 480855 44468 480869 44504
rect 480855 44457 480861 44468
rect 452399 44420 452405 44428
rect 452392 44384 452405 44420
rect 452399 44376 452405 44384
rect 452457 44420 452463 44428
rect 480881 44420 480887 44425
rect 452457 44384 480887 44420
rect 452457 44376 452463 44384
rect 480881 44373 480887 44384
rect 480939 44420 480945 44425
rect 480939 44384 480953 44420
rect 480939 44373 480945 44384
rect 447037 44336 447043 44344
rect 447019 44300 447043 44336
rect 447037 44292 447043 44300
rect 447095 44336 447101 44344
rect 480965 44336 480971 44341
rect 447095 44300 480971 44336
rect 447095 44292 447101 44300
rect 480965 44289 480971 44300
rect 481023 44336 481029 44341
rect 481023 44300 481037 44336
rect 481023 44289 481029 44300
rect 452237 44252 452243 44260
rect 452235 44216 452243 44252
rect 452237 44208 452243 44216
rect 452295 44252 452301 44260
rect 481049 44252 481055 44257
rect 452295 44216 481055 44252
rect 452295 44208 452301 44216
rect 481049 44205 481055 44216
rect 481107 44252 481113 44257
rect 481107 44216 481121 44252
rect 481107 44205 481113 44216
rect 447201 44168 447207 44176
rect 447177 44132 447207 44168
rect 447201 44124 447207 44132
rect 447259 44168 447265 44176
rect 481133 44168 481139 44173
rect 447259 44132 481139 44168
rect 447259 44124 447265 44132
rect 481133 44121 481139 44132
rect 481191 44168 481197 44173
rect 481191 44132 481205 44168
rect 481191 44121 481197 44132
rect 452082 44084 452088 44092
rect 452080 44048 452088 44084
rect 452082 44040 452088 44048
rect 452140 44084 452146 44092
rect 481217 44084 481223 44089
rect 452140 44048 481223 44084
rect 452140 44040 452146 44048
rect 481217 44037 481223 44048
rect 481275 44084 481281 44089
rect 481275 44048 481289 44084
rect 481275 44037 481281 44048
rect 447354 44000 447365 44008
rect 447345 43964 447365 44000
rect 447354 43956 447365 43964
rect 447417 44000 447423 44008
rect 481301 44000 481307 44005
rect 447417 43964 481307 44000
rect 447417 43956 447423 43964
rect 481301 43953 481307 43964
rect 481359 44000 481365 44005
rect 481359 43964 481373 44000
rect 481359 43953 481365 43964
rect 451914 43872 451920 43924
rect 451972 43916 451978 43924
rect 481385 43916 481391 43921
rect 451972 43880 481391 43916
rect 451972 43872 451978 43880
rect 481385 43869 481391 43880
rect 481443 43916 481449 43921
rect 481443 43880 481457 43916
rect 481443 43869 481449 43880
rect 447518 43832 447524 43840
rect 447507 43796 447524 43832
rect 447518 43788 447524 43796
rect 447576 43832 447582 43840
rect 481469 43832 481475 43837
rect 447576 43796 481475 43832
rect 447576 43788 447582 43796
rect 481469 43785 481475 43796
rect 481527 43832 481533 43837
rect 481527 43796 481541 43832
rect 481527 43785 481533 43796
rect 451759 43748 451765 43756
rect 451754 43712 451765 43748
rect 451759 43704 451765 43712
rect 451817 43748 451823 43756
rect 481553 43748 481559 43753
rect 451817 43712 481559 43748
rect 451817 43704 451823 43712
rect 481553 43701 481559 43712
rect 481611 43748 481617 43753
rect 481611 43712 481625 43748
rect 481611 43701 481617 43712
rect 447682 43664 447688 43672
rect 447664 43628 447688 43664
rect 447682 43620 447688 43628
rect 447740 43664 447746 43672
rect 481637 43664 481643 43669
rect 447740 43628 481643 43664
rect 447740 43620 447746 43628
rect 481637 43617 481643 43628
rect 481695 43664 481701 43669
rect 481695 43628 481709 43664
rect 481695 43617 481701 43628
rect 451597 43580 451603 43588
rect 451590 43544 451603 43580
rect 451597 43536 451603 43544
rect 451655 43580 451661 43588
rect 481721 43580 481727 43585
rect 451655 43544 481727 43580
rect 451655 43536 451661 43544
rect 481721 43533 481727 43544
rect 481779 43580 481785 43585
rect 481779 43544 481793 43580
rect 481779 43533 481785 43544
rect 447840 43496 447846 43504
rect 447819 43460 447846 43496
rect 447840 43452 447846 43460
rect 447898 43496 447904 43504
rect 481805 43496 481811 43501
rect 447898 43460 481811 43496
rect 447898 43452 447904 43460
rect 481805 43449 481811 43460
rect 481863 43449 481869 43501
rect 248253 42860 248259 42912
rect 248311 42904 248317 42912
rect 287758 42904 287764 42912
rect 248311 42868 255008 42904
rect 282220 42868 287764 42904
rect 248311 42860 248317 42868
rect 287758 42860 287764 42868
rect 287816 42860 287822 42912
rect 451969 42875 459639 43075
rect 248752 42776 248758 42828
rect 248810 42820 248816 42828
rect 288588 42820 288594 42828
rect 248810 42784 254993 42820
rect 282221 42784 288594 42820
rect 248810 42776 248816 42784
rect 288588 42776 288594 42784
rect 288646 42776 288652 42828
rect 249509 42692 249515 42744
rect 249567 42736 249573 42744
rect 289265 42736 289271 42744
rect 249567 42700 254970 42736
rect 282220 42700 289271 42736
rect 249567 42692 249573 42700
rect 289265 42692 289271 42700
rect 289323 42692 289329 42744
rect 353182 42652 353188 42660
rect 352466 42608 353188 42652
rect 353240 42608 353246 42660
rect 353266 42366 353272 42376
rect 352468 42324 353272 42366
rect 353324 42324 353330 42376
rect 352468 42320 353314 42324
rect 8350 41856 8356 41908
rect 8408 41896 8414 41908
rect 8408 41868 12964 41896
rect 8408 41856 8414 41868
rect 451969 41808 452125 42875
rect 459416 41808 459639 42875
rect 8462 41731 8468 41783
rect 8520 41771 8526 41783
rect 8520 41743 12967 41771
rect 8520 41731 8526 41743
rect 8574 41646 8580 41658
rect 8569 41618 8580 41646
rect 8574 41606 8580 41618
rect 8632 41646 8638 41658
rect 8632 41618 12970 41646
rect 8632 41606 8638 41618
rect 451969 41608 459639 41808
rect 472888 42852 480558 43008
rect 472888 41785 473111 42852
rect 480402 41785 480558 42852
rect 8686 41491 8692 41543
rect 8744 41531 8750 41543
rect 472888 41541 480558 41785
rect 541584 41605 541644 47124
rect 539822 41545 541644 41605
rect 541700 47052 568108 47058
rect 541700 47000 568048 47052
rect 568100 47000 568108 47052
rect 541700 46998 568108 47000
rect 8744 41503 12954 41531
rect 8744 41491 8750 41503
rect 541700 41485 541760 46998
rect 539834 41425 541760 41485
rect 567034 41424 567040 41436
rect 559906 41396 567040 41424
rect 567034 41384 567040 41396
rect 567092 41384 567098 41436
rect 567146 41302 567152 41314
rect 559892 41274 567152 41302
rect 567146 41262 567152 41274
rect 567204 41262 567210 41314
rect 566810 41170 566816 41182
rect 559896 41142 566816 41170
rect 566810 41130 566816 41142
rect 566868 41130 566874 41182
rect 566922 41066 566928 41078
rect 559916 41038 566928 41066
rect 566922 41026 566928 41038
rect 566980 41026 566986 41078
rect 83534 40578 83546 40630
rect 83598 40578 86019 40630
rect 353690 39418 353696 39426
rect 352502 39382 353696 39418
rect 353690 39374 353696 39382
rect 353748 39374 353754 39426
rect 353014 37670 353020 37682
rect 352468 37634 353020 37670
rect 353014 37630 353020 37634
rect 353072 37630 353078 37682
rect 353098 37380 353104 37394
rect 352474 37346 353104 37380
rect 353098 37342 353104 37346
rect 353156 37342 353162 37394
rect 7902 35945 7908 35997
rect 7960 35985 7966 35997
rect 7960 35957 12958 35985
rect 7960 35945 7966 35957
rect 8014 35824 8020 35876
rect 8072 35864 8078 35876
rect 8072 35836 12967 35864
rect 8072 35824 8078 35836
rect 8126 35706 8132 35758
rect 8184 35746 8190 35758
rect 8184 35718 12955 35746
rect 8184 35706 8190 35718
rect 539822 35639 543176 35699
rect 8238 35581 8244 35633
rect 8296 35621 8302 35633
rect 8296 35593 12974 35621
rect 8296 35581 8302 35593
rect 539814 35519 543072 35579
rect 543012 34620 543072 35519
rect 543116 34764 543176 35639
rect 566586 35518 566592 35530
rect 559868 35490 566592 35518
rect 566586 35478 566592 35490
rect 566644 35478 566650 35530
rect 566698 35390 566704 35402
rect 559918 35362 566704 35390
rect 566698 35350 566704 35362
rect 566756 35350 566762 35402
rect 566362 35284 566368 35296
rect 559930 35256 566368 35284
rect 566362 35244 566368 35256
rect 566420 35244 566426 35296
rect 566474 35144 566480 35156
rect 559930 35116 566480 35144
rect 566474 35104 566480 35116
rect 566532 35104 566538 35156
rect 543116 34756 568446 34764
rect 543116 34704 568384 34756
rect 568436 34704 568446 34756
rect 543012 34612 568556 34620
rect 543012 34560 568496 34612
rect 568548 34560 568556 34612
rect 353852 34422 353858 34430
rect 352376 34386 353858 34422
rect 353852 34378 353858 34386
rect 353910 34378 353916 34430
rect 542504 33520 568218 33528
rect 542504 33468 568160 33520
rect 568212 33468 568218 33520
rect 352846 32710 352852 32718
rect 352474 32666 352852 32710
rect 352904 32666 352910 32718
rect 352930 32418 352936 32428
rect 352468 32376 352936 32418
rect 352988 32376 352994 32428
rect 352468 32374 352978 32376
rect 273490 31314 273966 31318
rect 273478 31262 273484 31314
rect 273536 31262 273966 31314
rect 273490 31258 273966 31262
rect 273406 31193 273989 31198
rect 273394 31141 273400 31193
rect 273452 31141 273989 31193
rect 273406 31138 273989 31141
rect 353938 29476 353944 29484
rect 352350 29440 353944 29476
rect 353938 29432 353944 29440
rect 353996 29432 354002 29484
rect 233036 28376 233042 28384
rect 233034 28340 233042 28376
rect 233036 28332 233042 28340
rect 233094 28376 233100 28384
rect 233094 28340 234506 28376
rect 233094 28332 233100 28340
rect 173946 27872 173952 27924
rect 174004 27916 174010 27924
rect 177099 27916 177135 28103
rect 542504 28040 542564 33468
rect 539814 27980 542564 28040
rect 542634 33426 568330 33432
rect 542634 33374 568272 33426
rect 568324 33374 568330 33426
rect 542634 33372 568330 33374
rect 542634 27920 542694 33372
rect 566138 28026 566144 28038
rect 559632 27998 566144 28026
rect 566138 27986 566144 27998
rect 566196 27986 566202 28038
rect 174004 27880 177135 27916
rect 174004 27872 174010 27880
rect 539814 27860 542694 27920
rect 566250 27918 566256 27930
rect 559618 27890 566256 27918
rect 566250 27878 566256 27890
rect 566308 27878 566314 27930
rect 565914 27804 565920 27816
rect 559612 27776 565920 27804
rect 565914 27764 565920 27776
rect 565972 27764 565978 27816
rect 352678 27728 352684 27736
rect 7454 27666 7460 27718
rect 7512 27706 7518 27718
rect 7512 27678 12953 27706
rect 352470 27684 352684 27728
rect 352736 27684 352742 27736
rect 7512 27666 7518 27678
rect 566026 27674 566032 27686
rect 559584 27646 566032 27674
rect 566026 27634 566032 27646
rect 566084 27634 566090 27686
rect 7566 27540 7572 27592
rect 7624 27580 7630 27592
rect 7624 27552 12984 27580
rect 7624 27540 7630 27552
rect 7678 27413 7684 27465
rect 7736 27453 7742 27465
rect 7736 27425 12976 27453
rect 7736 27413 7742 27425
rect 352762 27424 352768 27432
rect 352470 27382 352768 27424
rect 352762 27380 352768 27382
rect 352820 27380 352826 27432
rect 7790 27290 7796 27342
rect 7848 27330 7854 27342
rect 7848 27302 12960 27330
rect 7848 27290 7854 27302
rect 257238 26004 257390 26022
rect 257238 24982 257258 26004
rect 257372 24982 257390 26004
rect 273656 25407 274016 25412
rect 273646 25355 273652 25407
rect 273704 25355 274016 25407
rect 273656 25352 274016 25355
rect 273574 25286 273966 25292
rect 273562 25234 273568 25286
rect 273620 25234 273966 25286
rect 273574 25232 273966 25234
rect 257238 24958 257390 24982
rect 354026 24522 354078 24528
rect 352416 24478 354026 24514
rect 354026 24464 354078 24470
rect 353518 22742 353524 22750
rect 352474 22698 353524 22742
rect 353576 22698 353582 22750
rect 431742 22602 439077 22807
rect 353602 22448 353608 22456
rect 352474 22406 353608 22448
rect 353602 22404 353608 22406
rect 353660 22404 353666 22456
rect 7230 21744 7236 21796
rect 7288 21784 7294 21796
rect 431742 21785 431923 22602
rect 438850 21785 439077 22602
rect 7288 21756 12981 21784
rect 7288 21744 7294 21756
rect 7342 21625 7348 21677
rect 7400 21665 7406 21677
rect 7400 21637 12986 21665
rect 7400 21625 7406 21637
rect 431742 21603 439077 21785
rect 472975 22662 478554 22814
rect 472975 21637 473177 22662
rect 478353 21637 478554 22662
rect 569274 22132 569280 22144
rect 539854 22088 540776 22116
rect 559602 22104 569280 22132
rect 569274 22092 569280 22104
rect 569332 22092 569338 22144
rect 539860 21970 540694 21998
rect 7006 21512 7012 21564
rect 7064 21552 7070 21564
rect 7064 21524 13080 21552
rect 7064 21512 7070 21524
rect 472975 21503 478554 21637
rect 540666 21550 540694 21970
rect 540748 21658 540776 22088
rect 569386 22010 569392 22022
rect 559578 21982 569392 22010
rect 569386 21970 569392 21982
rect 569444 21970 569450 22022
rect 568826 21878 568832 21890
rect 559620 21850 568832 21878
rect 568826 21838 568832 21850
rect 568884 21838 568890 21890
rect 568938 21776 568944 21788
rect 559606 21748 568944 21776
rect 568938 21736 568944 21748
rect 568996 21736 569002 21788
rect 569050 21658 569056 21670
rect 540748 21630 569056 21658
rect 569050 21618 569056 21630
rect 569108 21618 569114 21670
rect 569162 21550 569168 21562
rect 540666 21522 569168 21550
rect 569162 21510 569168 21522
rect 569220 21510 569226 21562
rect 7118 21391 7124 21443
rect 7176 21431 7182 21443
rect 7176 21403 13012 21431
rect 7176 21391 7182 21403
rect 530446 21341 530452 21349
rect 530443 21305 530452 21341
rect 467474 21290 467480 21299
rect 467468 21254 467480 21290
rect 467474 21247 467480 21254
rect 467532 21290 467538 21299
rect 530446 21297 530452 21305
rect 530504 21341 530510 21349
rect 540937 21341 540943 21349
rect 530504 21305 540943 21341
rect 530504 21297 530510 21305
rect 540937 21297 540943 21305
rect 540995 21341 541001 21349
rect 540995 21305 541009 21341
rect 540995 21297 541001 21305
rect 467532 21254 483856 21290
rect 530530 21257 530536 21265
rect 467532 21247 467538 21254
rect 465392 21206 465398 21213
rect 465386 21170 465398 21206
rect 465392 21161 465398 21170
rect 465450 21206 465456 21213
rect 465450 21170 483772 21206
rect 465450 21161 465456 21170
rect 465060 21122 465066 21128
rect 465053 21086 465066 21122
rect 465060 21076 465066 21086
rect 465118 21122 465124 21128
rect 465118 21086 483688 21122
rect 465118 21076 465124 21086
rect 464764 21038 464770 21047
rect 464758 21002 464770 21038
rect 464764 20995 464770 21002
rect 464822 21038 464828 21047
rect 464822 21002 483604 21038
rect 464822 20995 464828 21002
rect 464463 20954 464469 20961
rect 464455 20918 464469 20954
rect 464463 20909 464469 20918
rect 464521 20954 464527 20961
rect 464521 20918 483520 20954
rect 464521 20909 464527 20918
rect 482490 19988 482496 19996
rect 395426 19952 482496 19988
rect 354104 19610 354110 19618
rect 352458 19574 354110 19610
rect 354104 19566 354110 19574
rect 354162 19566 354168 19618
rect 354194 19498 354246 19504
rect 354188 19490 354194 19498
rect 352444 19454 354194 19490
rect 354188 19446 354194 19454
rect 354246 19446 354252 19498
rect 354194 19440 354246 19446
rect 354358 19304 354364 19356
rect 354416 19348 354422 19356
rect 395426 19348 395462 19952
rect 482490 19944 482496 19952
rect 482548 19944 482554 19996
rect 482406 19904 482412 19912
rect 354416 19312 395462 19348
rect 395510 19868 482412 19904
rect 354416 19304 354422 19312
rect 354274 19220 354280 19272
rect 354332 19264 354338 19272
rect 395510 19264 395546 19868
rect 482406 19860 482412 19868
rect 482464 19904 482470 19912
rect 482464 19868 482480 19904
rect 482464 19860 482470 19868
rect 482322 19820 482328 19828
rect 354332 19228 395546 19264
rect 395594 19784 482328 19820
rect 354332 19220 354338 19228
rect 294461 19081 295062 19197
rect 354190 19136 354196 19188
rect 354248 19180 354254 19188
rect 395594 19180 395630 19784
rect 482322 19776 482328 19784
rect 482380 19820 482386 19828
rect 482380 19784 482396 19820
rect 482380 19776 482386 19784
rect 482238 19736 482244 19744
rect 354248 19144 395630 19180
rect 395678 19700 482244 19736
rect 354248 19136 354254 19144
rect 294461 16433 294545 19081
rect 295010 16433 295062 19081
rect 354106 19052 354112 19104
rect 354164 19096 354170 19104
rect 395678 19096 395714 19700
rect 482238 19692 482244 19700
rect 482296 19736 482302 19744
rect 482296 19700 482312 19736
rect 482296 19692 482302 19700
rect 482154 19652 482160 19660
rect 354164 19060 395714 19096
rect 395762 19616 482160 19652
rect 354164 19052 354170 19060
rect 354022 18968 354028 19020
rect 354080 19012 354086 19020
rect 395762 19012 395798 19616
rect 482154 19608 482160 19616
rect 482212 19652 482218 19660
rect 482212 19616 482228 19652
rect 482212 19608 482218 19616
rect 482070 19568 482076 19576
rect 354080 18976 395798 19012
rect 395846 19532 482076 19568
rect 354080 18968 354086 18976
rect 353938 18884 353944 18936
rect 353996 18928 354002 18936
rect 395846 18928 395882 19532
rect 482070 19524 482076 19532
rect 482128 19568 482134 19576
rect 482128 19532 482144 19568
rect 482128 19524 482134 19532
rect 481986 19484 481992 19492
rect 353996 18892 395882 18928
rect 395930 19448 481992 19484
rect 353996 18884 354002 18892
rect 353854 18800 353860 18852
rect 353912 18844 353918 18852
rect 395930 18844 395966 19448
rect 481986 19440 481992 19448
rect 482044 19484 482050 19492
rect 482044 19448 482060 19484
rect 482044 19440 482050 19448
rect 481902 19400 481908 19408
rect 353912 18808 395966 18844
rect 396014 19364 481908 19400
rect 353912 18800 353918 18808
rect 353770 18716 353776 18768
rect 353828 18760 353834 18768
rect 396014 18760 396050 19364
rect 481902 19356 481908 19364
rect 481960 19400 481966 19408
rect 481960 19364 481976 19400
rect 481960 19356 481966 19364
rect 481818 19316 481824 19324
rect 353828 18724 396050 18760
rect 396098 19280 481824 19316
rect 353828 18716 353834 18724
rect 353686 18632 353692 18684
rect 353744 18676 353750 18684
rect 396098 18676 396134 19280
rect 481818 19272 481824 19280
rect 481876 19316 481882 19324
rect 481876 19280 481892 19316
rect 481876 19272 481882 19280
rect 481734 19232 481740 19240
rect 353744 18640 396134 18676
rect 396182 19196 481740 19232
rect 353744 18632 353750 18640
rect 353602 18548 353608 18600
rect 353660 18592 353666 18600
rect 396182 18592 396218 19196
rect 481734 19188 481740 19196
rect 481792 19232 481798 19240
rect 481792 19196 481808 19232
rect 481792 19188 481798 19196
rect 481650 19148 481656 19156
rect 353660 18556 396218 18592
rect 396266 19112 481656 19148
rect 353660 18548 353666 18556
rect 353518 18464 353524 18516
rect 353576 18508 353582 18516
rect 396266 18508 396302 19112
rect 481650 19104 481656 19112
rect 481708 19148 481714 19156
rect 481708 19112 481724 19148
rect 481708 19104 481714 19112
rect 481566 19064 481572 19072
rect 353576 18472 396302 18508
rect 396350 19028 481572 19064
rect 353576 18464 353582 18472
rect 353386 18380 353392 18432
rect 353444 18424 353450 18432
rect 396350 18424 396386 19028
rect 481566 19020 481572 19028
rect 481624 19064 481630 19072
rect 481624 19028 481640 19064
rect 481624 19020 481630 19028
rect 481482 18980 481488 18988
rect 353444 18388 396386 18424
rect 396434 18944 481488 18980
rect 353444 18380 353450 18388
rect 352566 18296 352572 18348
rect 352624 18340 352630 18348
rect 396434 18340 396470 18944
rect 481482 18936 481488 18944
rect 481540 18980 481546 18988
rect 481540 18944 481556 18980
rect 481540 18936 481546 18944
rect 481398 18896 481404 18904
rect 352624 18304 396470 18340
rect 396518 18860 481404 18896
rect 352624 18296 352630 18304
rect 353266 18212 353272 18264
rect 353324 18256 353330 18264
rect 396518 18256 396554 18860
rect 481398 18852 481404 18860
rect 481456 18896 481462 18904
rect 481456 18860 481472 18896
rect 481456 18852 481462 18860
rect 481314 18812 481320 18820
rect 353324 18220 396554 18256
rect 396602 18776 481320 18812
rect 353324 18212 353330 18220
rect 353182 18128 353188 18180
rect 353240 18172 353246 18180
rect 396602 18172 396638 18776
rect 481314 18768 481320 18776
rect 481372 18812 481378 18820
rect 481372 18776 481388 18812
rect 481372 18768 481378 18776
rect 481230 18728 481236 18736
rect 353240 18136 396638 18172
rect 396686 18692 481236 18728
rect 353240 18128 353246 18136
rect 353098 18044 353104 18096
rect 353156 18088 353162 18096
rect 396686 18088 396722 18692
rect 481230 18684 481236 18692
rect 481288 18728 481294 18736
rect 481288 18692 481304 18728
rect 481288 18684 481294 18692
rect 481146 18644 481152 18652
rect 353156 18052 396722 18088
rect 396770 18608 481152 18644
rect 353156 18044 353162 18052
rect 353014 17960 353020 18012
rect 353072 18004 353078 18012
rect 396770 18004 396806 18608
rect 481146 18600 481152 18608
rect 481204 18644 481210 18652
rect 481204 18608 481220 18644
rect 481204 18600 481210 18608
rect 481062 18560 481068 18568
rect 353072 17968 396806 18004
rect 396854 18524 481068 18560
rect 353072 17960 353078 17968
rect 352930 17876 352936 17928
rect 352988 17920 352994 17928
rect 396854 17920 396890 18524
rect 481062 18516 481068 18524
rect 481120 18560 481126 18568
rect 481120 18524 481136 18560
rect 481120 18516 481126 18524
rect 480978 18476 480984 18484
rect 352988 17884 396890 17920
rect 396938 18440 480984 18476
rect 352988 17876 352994 17884
rect 352846 17792 352852 17844
rect 352904 17836 352910 17844
rect 396938 17836 396974 18440
rect 480978 18432 480984 18440
rect 481036 18476 481042 18484
rect 481036 18440 481052 18476
rect 481036 18432 481042 18440
rect 480894 18392 480900 18400
rect 352904 17800 396974 17836
rect 397022 18356 480900 18392
rect 352904 17792 352910 17800
rect 352566 17776 352572 17784
rect 352466 17740 352572 17776
rect 352566 17732 352572 17740
rect 352624 17732 352630 17784
rect 352762 17708 352768 17760
rect 352820 17752 352826 17760
rect 397022 17752 397058 18356
rect 480894 18348 480900 18356
rect 480952 18392 480958 18400
rect 480952 18356 480968 18392
rect 480952 18348 480958 18356
rect 480810 18308 480816 18316
rect 352820 17716 397058 17752
rect 397106 18272 480816 18308
rect 352820 17708 352826 17716
rect 352678 17624 352684 17676
rect 352736 17668 352742 17676
rect 397106 17668 397142 18272
rect 480810 18264 480816 18272
rect 480868 18308 480874 18316
rect 480868 18272 480884 18308
rect 480868 18264 480874 18272
rect 352736 17632 397142 17668
rect 352736 17624 352742 17632
rect 353386 17496 353392 17504
rect 352458 17460 353392 17496
rect 353386 17452 353392 17460
rect 353444 17452 353450 17504
rect 294461 16310 295062 16433
rect 12607 16017 12613 16069
rect 12665 16062 12671 16069
rect 31206 16062 31212 16072
rect 12665 16026 31212 16062
rect 12665 16017 12671 16026
rect 31206 16020 31212 16026
rect 31264 16020 31270 16072
rect 12719 15933 12725 15985
rect 12777 15978 12783 15985
rect 31290 15978 31296 15988
rect 12777 15942 31296 15978
rect 12777 15933 12783 15942
rect 31290 15936 31296 15942
rect 31348 15936 31354 15988
rect 12831 15894 12837 15901
rect 12828 15858 12837 15894
rect 12831 15849 12837 15858
rect 12889 15894 12895 15901
rect 31374 15894 31380 15904
rect 12889 15858 31380 15894
rect 12889 15849 12895 15858
rect 31374 15852 31380 15858
rect 31432 15852 31438 15904
rect 12943 15765 12949 15817
rect 13001 15810 13007 15817
rect 31458 15810 31464 15820
rect 13001 15774 31464 15810
rect 13001 15765 13007 15774
rect 31458 15768 31464 15774
rect 31516 15768 31522 15820
rect 13055 15681 13061 15733
rect 13113 15726 13119 15733
rect 31542 15726 31548 15736
rect 13113 15690 31548 15726
rect 13113 15681 13119 15690
rect 31542 15684 31548 15690
rect 31600 15726 31606 15736
rect 367939 15732 367945 15849
rect 368062 15732 368068 15849
rect 31600 15690 31610 15726
rect 31600 15684 31606 15690
rect 13167 15597 13173 15649
rect 13225 15642 13231 15649
rect 31626 15642 31632 15652
rect 13225 15606 31632 15642
rect 13225 15597 13231 15606
rect 31626 15600 31632 15606
rect 31684 15642 31690 15652
rect 31684 15606 31694 15642
rect 31684 15600 31690 15606
rect 13954 15558 13960 15561
rect 13950 15522 13960 15558
rect 13954 15509 13960 15522
rect 14012 15558 14018 15561
rect 31710 15558 31716 15568
rect 14012 15522 31716 15558
rect 14012 15509 14018 15522
rect 31710 15516 31716 15522
rect 31768 15516 31774 15568
rect 14066 15425 14072 15477
rect 14124 15474 14130 15477
rect 31794 15474 31800 15484
rect 14124 15438 31800 15474
rect 14124 15425 14130 15438
rect 31794 15432 31800 15438
rect 31852 15432 31858 15484
rect 14178 15390 14184 15393
rect 14168 15354 14184 15390
rect 14178 15341 14184 15354
rect 14236 15390 14242 15393
rect 31878 15390 31884 15400
rect 14236 15354 31884 15390
rect 14236 15341 14242 15354
rect 31878 15348 31884 15354
rect 31936 15348 31942 15400
rect 14290 15306 14296 15309
rect 14288 15270 14296 15306
rect 14290 15257 14296 15270
rect 14348 15306 14354 15309
rect 31962 15306 31968 15316
rect 14348 15270 31968 15306
rect 14348 15257 14354 15270
rect 31962 15264 31968 15270
rect 32020 15264 32026 15316
rect 14402 15222 14408 15225
rect 14398 15186 14408 15222
rect 14402 15173 14408 15186
rect 14460 15222 14466 15225
rect 32046 15222 32052 15232
rect 14460 15186 32052 15222
rect 14460 15173 14466 15186
rect 32046 15180 32052 15186
rect 32104 15180 32110 15232
rect 14514 15138 14520 15141
rect 14510 15102 14520 15138
rect 14514 15089 14520 15102
rect 14572 15138 14578 15141
rect 32130 15138 32136 15148
rect 14572 15102 32136 15138
rect 14572 15089 14578 15102
rect 32130 15096 32136 15102
rect 32188 15096 32194 15148
rect 14626 15005 14632 15057
rect 14684 15054 14690 15057
rect 32214 15054 32220 15064
rect 14684 15018 32220 15054
rect 14684 15005 14690 15018
rect 32214 15012 32220 15018
rect 32272 15012 32278 15064
rect 14738 14970 14744 14973
rect 14732 14934 14744 14970
rect 14738 14921 14744 14934
rect 14796 14970 14802 14973
rect 32298 14970 32304 14980
rect 14796 14934 32304 14970
rect 14796 14921 14802 14934
rect 32298 14928 32304 14934
rect 32356 14928 32362 14980
rect 14850 14837 14856 14889
rect 14908 14886 14914 14889
rect 32382 14886 32388 14896
rect 14908 14850 32388 14886
rect 14908 14837 14914 14850
rect 32382 14844 32388 14850
rect 32440 14844 32446 14896
rect 14962 14802 14968 14805
rect 14958 14766 14968 14802
rect 14962 14753 14968 14766
rect 15020 14802 15026 14805
rect 32466 14802 32472 14812
rect 15020 14766 32472 14802
rect 15020 14753 15026 14766
rect 32466 14760 32472 14766
rect 32524 14760 32530 14812
rect 15073 14718 15079 14721
rect 15072 14682 15079 14718
rect 15073 14669 15079 14682
rect 15131 14718 15137 14721
rect 32550 14718 32556 14728
rect 15131 14682 32556 14718
rect 15131 14669 15137 14682
rect 32550 14676 32556 14682
rect 32608 14676 32614 14728
rect 15184 14585 15190 14637
rect 15242 14634 15248 14637
rect 32634 14634 32640 14644
rect 15242 14598 32640 14634
rect 15242 14585 15248 14598
rect 32634 14592 32640 14598
rect 32692 14592 32698 14644
rect 15295 14550 15301 14553
rect 15290 14514 15301 14550
rect 15295 14501 15301 14514
rect 15353 14550 15359 14553
rect 32718 14550 32724 14560
rect 15353 14514 32724 14550
rect 15353 14501 15359 14514
rect 32718 14508 32724 14514
rect 32776 14508 32782 14560
rect 15406 14466 15412 14469
rect 15404 14430 15412 14466
rect 15406 14417 15412 14430
rect 15464 14466 15470 14469
rect 32802 14466 32808 14476
rect 15464 14430 32808 14466
rect 15464 14417 15470 14430
rect 32802 14424 32808 14430
rect 32860 14466 32866 14476
rect 32860 14430 32868 14466
rect 32860 14424 32866 14430
rect 15517 14333 15523 14385
rect 15575 14382 15581 14385
rect 32886 14382 32892 14392
rect 15575 14346 32892 14382
rect 15575 14333 15581 14346
rect 32886 14340 32892 14346
rect 32944 14340 32950 14392
rect 15628 14249 15634 14301
rect 15686 14298 15692 14301
rect 32970 14298 32976 14308
rect 15686 14262 32976 14298
rect 15686 14249 15692 14262
rect 32970 14256 32976 14262
rect 33028 14256 33034 14308
rect 15739 14214 15745 14217
rect 15738 14178 15745 14214
rect 15739 14165 15745 14178
rect 15797 14214 15803 14217
rect 33054 14214 33060 14224
rect 15797 14178 33060 14214
rect 15797 14165 15803 14178
rect 33054 14172 33060 14178
rect 33112 14172 33118 14224
rect 15850 14130 15856 14133
rect 15844 14094 15856 14130
rect 15850 14081 15856 14094
rect 15908 14130 15914 14133
rect 33138 14130 33144 14140
rect 15908 14094 33144 14130
rect 15908 14081 15914 14094
rect 33138 14088 33144 14094
rect 33196 14088 33202 14140
rect 16198 14046 16204 14050
rect 16180 14010 16204 14046
rect 16198 13998 16204 14010
rect 16256 14046 16262 14050
rect 33222 14046 33228 14056
rect 16256 14010 33228 14046
rect 16256 13998 16262 14010
rect 33222 14004 33228 14010
rect 33280 14004 33286 14056
rect 16309 13962 16315 13966
rect 16304 13926 16315 13962
rect 16309 13914 16315 13926
rect 16367 13962 16373 13966
rect 33306 13962 33312 13972
rect 16367 13926 33312 13962
rect 16367 13914 16373 13926
rect 33306 13920 33312 13926
rect 33364 13920 33370 13972
rect 16420 13878 16426 13882
rect 16406 13842 16426 13878
rect 16420 13830 16426 13842
rect 16478 13878 16484 13882
rect 33390 13878 33396 13888
rect 16478 13842 33396 13878
rect 16478 13830 16484 13842
rect 33390 13836 33396 13842
rect 33448 13836 33454 13888
rect 16531 13794 16537 13798
rect 16522 13758 16537 13794
rect 16531 13746 16537 13758
rect 16589 13794 16595 13798
rect 33474 13794 33480 13804
rect 16589 13758 33480 13794
rect 16589 13746 16595 13758
rect 33474 13752 33480 13758
rect 33532 13752 33538 13804
rect 16642 13710 16648 13714
rect 16634 13674 16648 13710
rect 16642 13662 16648 13674
rect 16700 13710 16706 13714
rect 33558 13710 33564 13720
rect 16700 13674 33564 13710
rect 16700 13662 16706 13674
rect 33558 13668 33564 13674
rect 33616 13668 33622 13720
rect 16747 13586 16753 13638
rect 16805 13626 16811 13638
rect 33642 13626 33648 13636
rect 16805 13590 33648 13626
rect 16805 13586 16811 13590
rect 33642 13584 33648 13590
rect 33700 13584 33706 13636
rect 18878 13542 18884 13556
rect 18870 13506 18884 13542
rect 18878 13504 18884 13506
rect 18936 13542 18942 13556
rect 33726 13542 33732 13552
rect 18936 13506 33732 13542
rect 18936 13504 18942 13506
rect 33726 13500 33732 13506
rect 33784 13500 33790 13552
rect 363188 13493 363194 13545
rect 363246 13538 363252 13545
rect 363246 13499 363587 13538
rect 363246 13493 363252 13499
rect 18323 13458 18329 13466
rect 18314 13422 18329 13458
rect 18323 13414 18329 13422
rect 18381 13458 18387 13466
rect 33810 13458 33816 13468
rect 18381 13422 33816 13458
rect 18381 13414 18387 13422
rect 33810 13416 33816 13422
rect 33868 13416 33874 13468
rect 18434 13330 18440 13382
rect 18492 13374 18498 13382
rect 33894 13374 33900 13384
rect 18492 13338 33900 13374
rect 18492 13330 18498 13338
rect 33894 13332 33900 13338
rect 33952 13332 33958 13384
rect 18545 13246 18551 13298
rect 18603 13290 18609 13298
rect 33978 13290 33984 13300
rect 18603 13254 33984 13290
rect 18603 13246 18609 13254
rect 33978 13248 33984 13254
rect 34036 13290 34042 13300
rect 34036 13254 34048 13290
rect 34036 13248 34042 13254
rect 18656 13162 18662 13214
rect 18714 13206 18720 13214
rect 34062 13206 34068 13216
rect 18714 13170 34068 13206
rect 18714 13162 18720 13170
rect 34062 13164 34068 13170
rect 34120 13164 34126 13216
rect 18767 13078 18773 13130
rect 18825 13122 18831 13130
rect 34146 13122 34152 13132
rect 18825 13086 34152 13122
rect 18825 13078 18831 13086
rect 34146 13080 34152 13086
rect 34204 13122 34210 13132
rect 34204 13086 34216 13122
rect 34204 13080 34210 13086
rect 28510 12958 28516 12970
rect 28509 12922 28516 12958
rect 28510 12918 28516 12922
rect 28568 12958 28574 12970
rect 81824 12958 81830 12966
rect 28568 12922 81830 12958
rect 28568 12918 28574 12922
rect 81824 12914 81830 12922
rect 81882 12914 81888 12966
rect 28622 12874 28628 12886
rect 28613 12838 28628 12874
rect 28622 12834 28628 12838
rect 28680 12874 28686 12886
rect 81908 12874 81914 12882
rect 28680 12838 81914 12874
rect 28680 12834 28686 12838
rect 81908 12830 81914 12838
rect 81966 12830 81972 12882
rect 28734 12790 28740 12802
rect 28727 12754 28740 12790
rect 28734 12750 28740 12754
rect 28792 12790 28798 12802
rect 81992 12790 81998 12798
rect 28792 12754 81998 12790
rect 28792 12750 28798 12754
rect 81992 12746 81998 12754
rect 82050 12746 82056 12798
rect 28846 12706 28852 12717
rect 28842 12670 28852 12706
rect 28846 12665 28852 12670
rect 28904 12706 28910 12717
rect 82076 12706 82082 12714
rect 28904 12670 82082 12706
rect 28904 12665 28910 12670
rect 82076 12662 82082 12670
rect 82134 12662 82140 12714
rect 28958 12622 28964 12634
rect 28954 12586 28964 12622
rect 28958 12582 28964 12586
rect 29016 12622 29022 12634
rect 82160 12622 82166 12630
rect 29016 12586 82166 12622
rect 29016 12582 29022 12586
rect 82160 12578 82166 12586
rect 82218 12578 82224 12630
rect 29070 12538 29076 12550
rect 29067 12502 29076 12538
rect 29070 12498 29076 12502
rect 29128 12538 29134 12550
rect 82244 12538 82250 12546
rect 29128 12502 82250 12538
rect 29128 12498 29134 12502
rect 82244 12494 82250 12502
rect 82302 12494 82308 12546
rect 29182 12454 29188 12465
rect 29177 12418 29188 12454
rect 29182 12413 29188 12418
rect 29240 12454 29246 12465
rect 82328 12454 82334 12462
rect 29240 12418 82334 12454
rect 29240 12413 29246 12418
rect 82328 12410 82334 12418
rect 82386 12410 82392 12462
rect 29294 12370 29300 12381
rect 29291 12334 29300 12370
rect 29294 12329 29300 12334
rect 29352 12370 29358 12381
rect 82412 12370 82418 12378
rect 29352 12334 82418 12370
rect 29352 12329 29358 12334
rect 82412 12326 82418 12334
rect 82470 12326 82476 12378
rect 28398 12286 28404 12297
rect 28397 12250 28404 12286
rect 28398 12245 28404 12250
rect 28456 12286 28462 12297
rect 82496 12286 82502 12294
rect 28456 12250 82502 12286
rect 28456 12245 28462 12250
rect 82496 12242 82502 12250
rect 82554 12242 82560 12294
rect 28286 12202 28292 12213
rect 28281 12166 28292 12202
rect 28286 12161 28292 12166
rect 28344 12202 28350 12213
rect 82580 12202 82586 12210
rect 28344 12166 82586 12202
rect 28344 12161 28350 12166
rect 82580 12158 82586 12166
rect 82638 12158 82644 12210
rect 28174 12118 28180 12130
rect 28167 12082 28180 12118
rect 28174 12078 28180 12082
rect 28232 12118 28238 12130
rect 82664 12118 82670 12126
rect 28232 12082 82670 12118
rect 28232 12078 28238 12082
rect 82664 12074 82670 12082
rect 82722 12074 82728 12126
rect 28062 12034 28068 12045
rect 28058 11998 28068 12034
rect 28062 11993 28068 11998
rect 28120 12034 28126 12045
rect 82748 12034 82754 12042
rect 28120 11998 82754 12034
rect 28120 11993 28126 11998
rect 82748 11990 82754 11998
rect 82806 11990 82812 12042
rect 27950 11950 27956 11962
rect 27945 11914 27956 11950
rect 27950 11910 27956 11914
rect 28008 11950 28014 11962
rect 82832 11950 82838 11958
rect 28008 11914 82838 11950
rect 28008 11910 28014 11914
rect 82832 11906 82838 11914
rect 82890 11906 82896 11958
rect 27838 11866 27844 11880
rect 27833 11830 27844 11866
rect 27838 11828 27844 11830
rect 27896 11866 27902 11880
rect 82916 11866 82922 11874
rect 27896 11830 82922 11866
rect 27896 11828 27902 11830
rect 82916 11822 82922 11830
rect 82974 11822 82980 11874
rect 363274 11863 363280 11915
rect 363332 11910 363338 11915
rect 363332 11867 363583 11910
rect 363332 11863 363338 11867
rect 27726 11782 27732 11793
rect 27720 11746 27732 11782
rect 27726 11741 27732 11746
rect 27784 11782 27790 11793
rect 83000 11782 83006 11790
rect 27784 11746 83006 11782
rect 27784 11741 27790 11746
rect 83000 11738 83006 11746
rect 83058 11738 83064 11790
rect 27614 11658 27620 11710
rect 27672 11698 27678 11710
rect 83084 11698 83090 11706
rect 27672 11662 83090 11698
rect 27672 11658 27678 11662
rect 83084 11654 83090 11662
rect 83142 11654 83148 11706
rect 29851 11622 29857 11630
rect 29847 11586 29857 11622
rect 29851 11578 29857 11586
rect 29909 11622 29915 11630
rect 80943 11622 80949 11630
rect 29909 11587 80949 11622
rect 29909 11586 30629 11587
rect 30714 11586 80949 11587
rect 29909 11578 29915 11586
rect 80943 11578 80949 11586
rect 81001 11622 81007 11630
rect 81001 11586 81010 11622
rect 81001 11578 81007 11586
rect 30640 11538 30646 11546
rect 30632 11502 30646 11538
rect 30640 11494 30646 11502
rect 30698 11538 30704 11546
rect 81027 11538 81033 11546
rect 30698 11502 81033 11538
rect 30698 11494 30704 11502
rect 81027 11494 81033 11502
rect 81085 11538 81091 11546
rect 81085 11502 81094 11538
rect 81085 11494 81091 11502
rect 30526 11454 30532 11462
rect 30520 11418 30532 11454
rect 30526 11410 30532 11418
rect 30584 11454 30590 11462
rect 81111 11454 81117 11462
rect 30584 11418 81117 11454
rect 30584 11410 30590 11418
rect 81111 11410 81117 11418
rect 81169 11454 81175 11462
rect 81169 11418 81178 11454
rect 81169 11410 81175 11418
rect 30302 11370 30308 11378
rect 30297 11334 30308 11370
rect 30302 11326 30308 11334
rect 30360 11370 30366 11378
rect 81195 11370 81201 11378
rect 30360 11334 81201 11370
rect 30360 11326 30366 11334
rect 81195 11326 81201 11334
rect 81253 11370 81259 11378
rect 81253 11334 81262 11370
rect 81253 11326 81259 11334
rect 30411 11286 30417 11294
rect 30408 11250 30417 11286
rect 30411 11242 30417 11250
rect 30469 11286 30475 11294
rect 81279 11286 81285 11294
rect 30469 11250 81285 11286
rect 30469 11242 30475 11250
rect 81279 11242 81285 11250
rect 81337 11286 81343 11294
rect 81337 11250 81346 11286
rect 81337 11242 81343 11250
rect 30972 11202 30978 11210
rect 30967 11166 30978 11202
rect 30972 11158 30978 11166
rect 31030 11202 31036 11210
rect 81363 11202 81369 11210
rect 31030 11166 81369 11202
rect 31030 11158 31036 11166
rect 81363 11158 81369 11166
rect 81421 11202 81427 11210
rect 81421 11166 81430 11202
rect 81421 11158 81427 11166
rect 30863 11118 30869 11126
rect 30860 11082 30869 11118
rect 30863 11074 30869 11082
rect 30921 11118 30927 11126
rect 81447 11118 81453 11126
rect 30921 11082 81453 11118
rect 30921 11074 30927 11082
rect 81447 11074 81453 11082
rect 81505 11118 81511 11126
rect 81505 11082 81514 11118
rect 81505 11074 81511 11082
rect 31424 11034 31430 11042
rect 31421 10998 31430 11034
rect 31424 10990 31430 10998
rect 31482 11034 31488 11042
rect 81531 11034 81537 11042
rect 31482 10998 81537 11034
rect 31482 10990 31488 10998
rect 81531 10990 81537 10998
rect 81589 11034 81595 11042
rect 81589 10998 81598 11034
rect 81589 10990 81595 10998
rect 93473 10982 93509 11006
rect 95101 10982 95137 11006
rect 96729 10982 96765 11006
rect 98357 10982 98393 11006
rect 99985 10982 100021 11006
rect 101613 10982 101649 11006
rect 103241 10982 103277 11006
rect 104869 10982 104905 11006
rect 110099 10986 110174 10996
rect 30750 10950 30756 10958
rect 30746 10914 30756 10950
rect 30750 10906 30756 10914
rect 30808 10950 30814 10958
rect 81615 10950 81621 10958
rect 30808 10914 81621 10950
rect 30808 10906 30814 10914
rect 81615 10906 81621 10914
rect 81673 10950 81679 10958
rect 81673 10914 81682 10950
rect 92022 10930 92028 10982
rect 92080 10930 92086 10982
rect 93460 10930 93466 10982
rect 93518 10930 93524 10982
rect 95088 10930 95094 10982
rect 95146 10930 95152 10982
rect 96716 10930 96722 10982
rect 96774 10930 96780 10982
rect 98344 10930 98350 10982
rect 98402 10930 98408 10982
rect 99972 10930 99978 10982
rect 100030 10930 100036 10982
rect 101600 10930 101606 10982
rect 101658 10930 101664 10982
rect 103228 10930 103234 10982
rect 103286 10930 103292 10982
rect 104856 10930 104862 10982
rect 104914 10930 104920 10982
rect 93473 10928 93509 10930
rect 95101 10928 95137 10930
rect 96729 10928 96765 10930
rect 98357 10928 98393 10930
rect 99985 10928 100021 10930
rect 101613 10928 101649 10930
rect 103241 10928 103277 10930
rect 104869 10928 104905 10930
rect 110099 10928 110109 10986
rect 110167 10928 110174 10986
rect 110099 10921 110174 10928
rect 111727 10986 111802 10996
rect 111727 10928 111737 10986
rect 111795 10928 111802 10986
rect 111727 10921 111802 10928
rect 113355 10986 113430 10996
rect 113355 10928 113365 10986
rect 113423 10928 113430 10986
rect 113355 10921 113430 10928
rect 114983 10986 115058 10996
rect 114983 10928 114993 10986
rect 115051 10928 115058 10986
rect 114983 10921 115058 10928
rect 116611 10986 116686 10996
rect 116611 10928 116621 10986
rect 116679 10928 116686 10986
rect 116611 10921 116686 10928
rect 118239 10986 118314 10996
rect 118239 10928 118249 10986
rect 118307 10928 118314 10986
rect 118239 10921 118314 10928
rect 119867 10986 119942 10996
rect 119867 10928 119877 10986
rect 119935 10928 119942 10986
rect 119867 10921 119942 10928
rect 121494 10986 121569 10995
rect 121494 10928 121505 10986
rect 121563 10928 121569 10986
rect 121494 10920 121569 10928
rect 81673 10906 81679 10914
rect 31196 10866 31202 10874
rect 31190 10830 31202 10866
rect 31196 10822 31202 10830
rect 31254 10866 31260 10874
rect 81699 10866 81705 10874
rect 31254 10830 81705 10866
rect 31254 10822 31260 10830
rect 81699 10822 81705 10830
rect 81757 10866 81763 10874
rect 81757 10830 81766 10866
rect 81757 10822 81763 10830
rect 23022 10782 23028 10798
rect 23012 10746 23028 10782
rect 23080 10782 23086 10798
rect 122953 10782 122989 10973
rect 23080 10746 122989 10782
rect 23134 10698 23140 10707
rect 23132 10662 23140 10698
rect 23134 10655 23140 10662
rect 23192 10698 23198 10707
rect 23192 10662 122883 10698
rect 23192 10655 23198 10662
rect 23246 10614 23252 10626
rect 23244 10578 23252 10614
rect 23246 10574 23252 10578
rect 23304 10614 23310 10626
rect 23304 10578 122883 10614
rect 23304 10574 23310 10578
rect 23358 10530 23364 10545
rect 23356 10494 23364 10530
rect 23358 10493 23364 10494
rect 23416 10530 23422 10545
rect 23416 10494 122883 10530
rect 23416 10493 23422 10494
rect 23470 10446 23476 10456
rect 23468 10410 23476 10446
rect 23470 10404 23476 10410
rect 23528 10446 23534 10456
rect 23528 10410 122883 10446
rect 23528 10404 23534 10410
rect 23582 10362 23588 10373
rect 23580 10326 23588 10362
rect 23582 10321 23588 10326
rect 23640 10362 23646 10373
rect 121499 10362 121505 10377
rect 23640 10326 121505 10362
rect 23640 10321 23646 10326
rect 121499 10319 121505 10326
rect 121563 10362 121569 10377
rect 121563 10326 121571 10362
rect 121563 10319 121569 10326
rect 23694 10278 23700 10288
rect 23692 10242 23700 10278
rect 23694 10236 23700 10242
rect 23752 10278 23758 10288
rect 119871 10278 119877 10287
rect 23752 10242 119877 10278
rect 23752 10236 23758 10242
rect 119871 10229 119877 10242
rect 119935 10278 119941 10287
rect 119935 10242 119958 10278
rect 119935 10229 119941 10242
rect 23812 10204 23864 10210
rect 23804 10158 23812 10194
rect 118242 10194 118248 10207
rect 23864 10158 118248 10194
rect 118242 10155 118248 10158
rect 118300 10194 118306 10207
rect 118300 10158 118330 10194
rect 118300 10155 118306 10158
rect 23812 10146 23864 10152
rect 23924 10124 23976 10130
rect 23916 10074 23924 10110
rect 116614 10110 116620 10119
rect 23976 10074 116620 10110
rect 23924 10066 23976 10072
rect 116614 10067 116620 10074
rect 116672 10110 116678 10119
rect 116672 10074 116702 10110
rect 116672 10067 116678 10074
rect 24030 10026 24036 10041
rect 24028 9990 24036 10026
rect 24030 9989 24036 9990
rect 24088 10026 24094 10041
rect 114986 10026 114992 10040
rect 24088 9990 114992 10026
rect 24088 9989 24094 9990
rect 114986 9988 114992 9990
rect 115044 10026 115050 10040
rect 115044 9990 115074 10026
rect 115044 9988 115050 9990
rect 113364 9956 113416 9962
rect 24142 9942 24148 9956
rect 24140 9906 24148 9942
rect 24142 9904 24148 9906
rect 24200 9942 24206 9956
rect 24200 9906 113364 9942
rect 24200 9904 24206 9906
rect 113416 9906 113446 9942
rect 113364 9898 113416 9904
rect 24254 9858 24260 9870
rect 24252 9822 24260 9858
rect 24254 9818 24260 9822
rect 24312 9858 24318 9870
rect 111730 9858 111736 9870
rect 24312 9822 111736 9858
rect 24312 9818 24318 9822
rect 111730 9818 111736 9822
rect 111788 9858 111794 9870
rect 111788 9822 111818 9858
rect 111788 9818 111794 9822
rect 24366 9774 24372 9787
rect 24364 9738 24372 9774
rect 24366 9735 24372 9738
rect 24424 9774 24430 9787
rect 110102 9774 110108 9785
rect 24424 9738 110108 9774
rect 24424 9735 24430 9738
rect 110102 9733 110108 9738
rect 110160 9774 110166 9785
rect 110160 9738 110190 9774
rect 110160 9733 110166 9738
rect 24478 9690 24484 9702
rect 24476 9654 24484 9690
rect 24478 9650 24484 9654
rect 24536 9690 24542 9702
rect 92022 9690 92028 9698
rect 24536 9654 92028 9690
rect 24536 9650 24542 9654
rect 92022 9646 92028 9654
rect 92080 9690 92086 9698
rect 92080 9654 92094 9690
rect 92080 9646 92086 9654
rect 24590 9606 24596 9620
rect 24588 9570 24596 9606
rect 24590 9568 24596 9570
rect 24648 9606 24654 9620
rect 24648 9570 92184 9606
rect 24648 9568 24654 9570
rect 24702 9522 24708 9532
rect 24700 9486 24708 9522
rect 24702 9480 24708 9486
rect 24760 9522 24766 9532
rect 24760 9486 92184 9522
rect 24760 9480 24766 9486
rect 24814 9438 24820 9451
rect 24812 9402 24820 9438
rect 24814 9399 24820 9402
rect 24872 9438 24878 9451
rect 24872 9402 92184 9438
rect 24872 9399 24878 9402
rect 24926 9354 24932 9366
rect 24924 9318 24932 9354
rect 24926 9314 24932 9318
rect 24984 9354 24990 9366
rect 24984 9318 92184 9354
rect 24984 9314 24990 9318
rect 25038 9270 25044 9282
rect 25036 9234 25044 9270
rect 25038 9230 25044 9234
rect 25096 9270 25102 9282
rect 93460 9270 93466 9278
rect 25096 9234 93466 9270
rect 25096 9230 25102 9234
rect 93460 9226 93466 9234
rect 93518 9270 93524 9278
rect 93518 9234 93536 9270
rect 93518 9226 93524 9234
rect 25150 9186 25156 9198
rect 25148 9150 25156 9186
rect 25150 9146 25156 9150
rect 25208 9186 25214 9198
rect 95088 9186 95094 9195
rect 25208 9150 95094 9186
rect 25208 9146 25214 9150
rect 95088 9143 95094 9150
rect 95146 9186 95152 9195
rect 95146 9150 95186 9186
rect 95146 9143 95152 9150
rect 25262 9102 25268 9113
rect 25260 9066 25268 9102
rect 25262 9061 25268 9066
rect 25320 9102 25326 9113
rect 96716 9102 96722 9107
rect 25320 9066 96722 9102
rect 25320 9061 25326 9066
rect 96716 9055 96722 9066
rect 96774 9102 96780 9107
rect 96774 9066 96792 9102
rect 96774 9055 96780 9066
rect 483484 9033 483520 20918
rect 483568 9117 483604 21002
rect 483652 9201 483688 21086
rect 483736 9285 483772 21170
rect 483820 9369 483856 21254
rect 530527 21221 530536 21257
rect 530530 21213 530536 21221
rect 530588 21257 530594 21265
rect 541021 21257 541027 21265
rect 530588 21221 541027 21257
rect 530588 21213 530594 21221
rect 541021 21213 541027 21221
rect 541079 21257 541085 21265
rect 541079 21221 541093 21257
rect 541079 21213 541085 21221
rect 530614 21173 530620 21181
rect 530611 21137 530620 21173
rect 530614 21129 530620 21137
rect 530672 21173 530678 21181
rect 541105 21173 541111 21181
rect 530672 21137 541111 21173
rect 530672 21129 530678 21137
rect 541105 21129 541111 21137
rect 541163 21173 541169 21181
rect 541163 21137 541177 21173
rect 541163 21129 541169 21137
rect 530698 21089 530704 21097
rect 530695 21053 530704 21089
rect 530698 21045 530704 21053
rect 530756 21089 530762 21097
rect 541189 21089 541195 21097
rect 530756 21053 541195 21089
rect 530756 21045 530762 21053
rect 541189 21045 541195 21053
rect 541247 21089 541253 21097
rect 541247 21053 541261 21089
rect 541247 21045 541253 21053
rect 530782 21005 530788 21013
rect 530779 20969 530788 21005
rect 530782 20961 530788 20969
rect 530840 21005 530846 21013
rect 541273 21005 541279 21013
rect 530840 20969 541279 21005
rect 530840 20961 530846 20969
rect 541273 20961 541279 20969
rect 541331 21005 541337 21013
rect 541331 20969 541345 21005
rect 541331 20961 541337 20969
rect 530866 20921 530872 20929
rect 530863 20885 530872 20921
rect 530866 20877 530872 20885
rect 530924 20921 530930 20929
rect 541357 20921 541363 20929
rect 530924 20885 541363 20921
rect 530924 20877 530930 20885
rect 541357 20877 541363 20885
rect 541415 20921 541421 20929
rect 541415 20885 541429 20921
rect 541415 20877 541421 20885
rect 530950 20837 530956 20845
rect 530947 20801 530956 20837
rect 530950 20793 530956 20801
rect 531008 20837 531014 20845
rect 541441 20837 541447 20845
rect 531008 20801 541447 20837
rect 531008 20793 531014 20801
rect 541441 20793 541447 20801
rect 541499 20837 541505 20845
rect 541499 20801 541513 20837
rect 541499 20793 541505 20801
rect 531034 20753 531040 20761
rect 531031 20717 531040 20753
rect 531034 20709 531040 20717
rect 531092 20753 531098 20761
rect 541525 20753 541531 20761
rect 531092 20717 541531 20753
rect 531092 20709 531098 20717
rect 541525 20709 541531 20717
rect 541583 20753 541589 20761
rect 541583 20717 541597 20753
rect 541583 20709 541589 20717
rect 531118 20669 531124 20677
rect 531115 20633 531124 20669
rect 531118 20625 531124 20633
rect 531176 20669 531182 20677
rect 541609 20669 541615 20677
rect 531176 20633 541615 20669
rect 531176 20625 531182 20633
rect 541609 20625 541615 20633
rect 541667 20669 541673 20677
rect 541667 20633 541681 20669
rect 541667 20625 541673 20633
rect 531202 20585 531208 20593
rect 531199 20549 531208 20585
rect 531202 20541 531208 20549
rect 531260 20585 531266 20593
rect 541693 20585 541699 20593
rect 531260 20549 541699 20585
rect 531260 20541 531266 20549
rect 541693 20541 541699 20549
rect 541751 20585 541757 20593
rect 541751 20549 541765 20585
rect 541751 20541 541757 20549
rect 531286 20501 531292 20509
rect 531283 20465 531292 20501
rect 531286 20457 531292 20465
rect 531344 20501 531350 20509
rect 541777 20501 541783 20509
rect 531344 20465 541783 20501
rect 531344 20457 531350 20465
rect 541777 20457 541783 20465
rect 541835 20501 541841 20509
rect 541835 20465 541849 20501
rect 541835 20457 541841 20465
rect 531370 20417 531376 20425
rect 531367 20381 531376 20417
rect 531370 20373 531376 20381
rect 531428 20417 531434 20425
rect 541861 20417 541867 20425
rect 531428 20381 541867 20417
rect 531428 20373 531434 20381
rect 541861 20373 541867 20381
rect 541919 20417 541925 20425
rect 541919 20381 541933 20417
rect 541919 20373 541925 20381
rect 531454 20333 531460 20341
rect 531451 20297 531460 20333
rect 531454 20289 531460 20297
rect 531512 20333 531518 20341
rect 541945 20333 541951 20341
rect 531512 20297 541951 20333
rect 531512 20289 531518 20297
rect 541945 20289 541951 20297
rect 542003 20333 542009 20341
rect 542003 20297 542017 20333
rect 542003 20289 542009 20297
rect 531538 20249 531544 20257
rect 531535 20213 531544 20249
rect 531538 20205 531544 20213
rect 531596 20249 531602 20257
rect 542029 20249 542035 20257
rect 531596 20213 542035 20249
rect 531596 20205 531602 20213
rect 542029 20205 542035 20213
rect 542087 20249 542093 20257
rect 542087 20213 542101 20249
rect 542087 20205 542093 20213
rect 531622 20165 531628 20173
rect 531619 20129 531628 20165
rect 531622 20121 531628 20129
rect 531680 20165 531686 20173
rect 542113 20165 542119 20173
rect 531680 20129 542119 20165
rect 531680 20121 531686 20129
rect 542113 20121 542119 20129
rect 542171 20165 542177 20173
rect 542171 20129 542185 20165
rect 542171 20121 542177 20129
rect 531706 20081 531712 20089
rect 531703 20045 531712 20081
rect 531706 20037 531712 20045
rect 531764 20081 531770 20089
rect 542197 20081 542203 20089
rect 531764 20045 542203 20081
rect 531764 20037 531770 20045
rect 542197 20037 542203 20045
rect 542255 20081 542261 20089
rect 542255 20045 542269 20081
rect 542255 20037 542261 20045
rect 531790 19997 531796 20005
rect 531787 19961 531796 19997
rect 531790 19953 531796 19961
rect 531848 19997 531854 20005
rect 542281 19997 542287 20005
rect 531848 19961 542287 19997
rect 531848 19953 531854 19961
rect 542281 19953 542287 19961
rect 542339 19997 542345 20005
rect 542339 19961 542353 19997
rect 542339 19953 542345 19961
rect 531874 19913 531880 19921
rect 531871 19877 531880 19913
rect 531874 19869 531880 19877
rect 531932 19913 531938 19921
rect 542365 19913 542371 19921
rect 531932 19877 542371 19913
rect 531932 19869 531938 19877
rect 542365 19869 542371 19877
rect 542423 19913 542429 19921
rect 542423 19877 542437 19913
rect 542423 19869 542429 19877
rect 531958 19829 531964 19837
rect 531955 19793 531964 19829
rect 531958 19785 531964 19793
rect 532016 19829 532022 19837
rect 542449 19829 542455 19837
rect 532016 19793 542455 19829
rect 532016 19785 532022 19793
rect 542449 19785 542455 19793
rect 542507 19829 542513 19837
rect 542507 19793 542521 19829
rect 542507 19785 542513 19793
rect 532042 19745 532048 19753
rect 532039 19709 532048 19745
rect 532042 19701 532048 19709
rect 532100 19745 532106 19753
rect 542533 19745 542539 19753
rect 532100 19709 542539 19745
rect 532100 19701 532106 19709
rect 542533 19701 542539 19709
rect 542591 19745 542597 19753
rect 542591 19709 542605 19745
rect 542591 19701 542597 19709
rect 532126 19661 532132 19669
rect 532123 19625 532132 19661
rect 532126 19617 532132 19625
rect 532184 19661 532190 19669
rect 542617 19661 542623 19669
rect 532184 19625 542623 19661
rect 532184 19617 532190 19625
rect 542617 19617 542623 19625
rect 542675 19661 542681 19669
rect 542675 19625 542689 19661
rect 542675 19617 542681 19625
rect 532210 19577 532216 19585
rect 532207 19541 532216 19577
rect 532210 19533 532216 19541
rect 532268 19577 532274 19585
rect 542701 19577 542707 19585
rect 532268 19541 542707 19577
rect 532268 19533 532274 19541
rect 542701 19533 542707 19541
rect 542759 19577 542765 19585
rect 542759 19541 542773 19577
rect 542759 19533 542765 19541
rect 532294 19493 532300 19501
rect 532291 19457 532300 19493
rect 532294 19449 532300 19457
rect 532352 19493 532358 19501
rect 542785 19493 542791 19501
rect 532352 19457 542791 19493
rect 532352 19449 532358 19457
rect 542785 19449 542791 19457
rect 542843 19493 542849 19501
rect 542843 19457 542857 19493
rect 542843 19449 542849 19457
rect 532378 19409 532384 19417
rect 532375 19373 532384 19409
rect 532378 19365 532384 19373
rect 532436 19409 532442 19417
rect 542869 19409 542875 19417
rect 532436 19373 542875 19409
rect 532436 19365 532442 19373
rect 542869 19365 542875 19373
rect 542927 19409 542933 19417
rect 542927 19373 542941 19409
rect 542927 19365 542933 19373
rect 532462 19325 532468 19333
rect 532459 19289 532468 19325
rect 532462 19281 532468 19289
rect 532520 19325 532526 19333
rect 542953 19325 542959 19333
rect 532520 19289 542959 19325
rect 532520 19281 532526 19289
rect 542953 19281 542959 19289
rect 543011 19325 543017 19333
rect 543011 19289 543025 19325
rect 543011 19281 543017 19289
rect 532546 19241 532552 19249
rect 532543 19205 532552 19241
rect 532546 19197 532552 19205
rect 532604 19241 532610 19249
rect 543037 19241 543043 19249
rect 532604 19205 543043 19241
rect 532604 19197 532610 19205
rect 543037 19197 543043 19205
rect 543095 19241 543101 19249
rect 543095 19205 543109 19241
rect 543095 19197 543101 19205
rect 532630 19157 532636 19165
rect 532627 19121 532636 19157
rect 532630 19113 532636 19121
rect 532688 19157 532694 19165
rect 543121 19157 543127 19165
rect 532688 19121 543127 19157
rect 532688 19113 532694 19121
rect 543121 19113 543127 19121
rect 543179 19157 543185 19165
rect 543179 19121 543193 19157
rect 543179 19113 543185 19121
rect 532714 19073 532720 19081
rect 532711 19037 532720 19073
rect 532714 19029 532720 19037
rect 532772 19073 532778 19081
rect 543205 19073 543211 19081
rect 532772 19037 543211 19073
rect 532772 19029 532778 19037
rect 543205 19029 543211 19037
rect 543263 19073 543269 19081
rect 543263 19037 543277 19073
rect 543263 19029 543269 19037
rect 532798 18989 532804 18997
rect 532795 18953 532804 18989
rect 532798 18945 532804 18953
rect 532856 18989 532862 18997
rect 543289 18989 543295 18997
rect 532856 18953 543295 18989
rect 532856 18945 532862 18953
rect 543289 18945 543295 18953
rect 543347 18989 543353 18997
rect 543347 18953 543361 18989
rect 543347 18945 543353 18953
rect 532882 18905 532888 18913
rect 532879 18869 532888 18905
rect 532882 18861 532888 18869
rect 532940 18905 532946 18913
rect 543373 18905 543379 18913
rect 532940 18869 543379 18905
rect 532940 18861 532946 18869
rect 543373 18861 543379 18869
rect 543431 18905 543437 18913
rect 543431 18869 543445 18905
rect 543431 18861 543437 18869
rect 532966 18821 532972 18829
rect 532963 18785 532972 18821
rect 532966 18777 532972 18785
rect 533024 18821 533030 18829
rect 543457 18821 543463 18829
rect 533024 18785 543463 18821
rect 533024 18777 533030 18785
rect 543457 18777 543463 18785
rect 543515 18821 543521 18829
rect 543515 18785 543529 18821
rect 543515 18777 543521 18785
rect 533050 18737 533056 18745
rect 533047 18701 533056 18737
rect 533050 18693 533056 18701
rect 533108 18737 533114 18745
rect 543541 18737 543547 18745
rect 533108 18701 543547 18737
rect 533108 18693 533114 18701
rect 543541 18693 543547 18701
rect 543599 18737 543605 18745
rect 543599 18701 543613 18737
rect 543599 18693 543605 18701
rect 533134 18653 533140 18661
rect 533131 18617 533140 18653
rect 533134 18609 533140 18617
rect 533192 18653 533198 18661
rect 543625 18653 543631 18661
rect 533192 18617 543631 18653
rect 533192 18609 533198 18617
rect 543625 18609 543631 18617
rect 543683 18653 543689 18661
rect 543683 18617 543697 18653
rect 543683 18609 543689 18617
rect 533218 18569 533224 18577
rect 533215 18533 533224 18569
rect 533218 18525 533224 18533
rect 533276 18569 533282 18577
rect 543709 18569 543715 18577
rect 533276 18533 543715 18569
rect 533276 18525 533282 18533
rect 543709 18525 543715 18533
rect 543767 18569 543773 18577
rect 543767 18533 543781 18569
rect 543767 18525 543773 18533
rect 533302 18485 533308 18493
rect 533299 18449 533308 18485
rect 533302 18441 533308 18449
rect 533360 18485 533366 18493
rect 543793 18485 543799 18493
rect 533360 18449 543799 18485
rect 533360 18441 533366 18449
rect 543793 18441 543799 18449
rect 543851 18441 543857 18493
rect 530252 18359 530258 18367
rect 530250 18323 530258 18359
rect 530252 18315 530258 18323
rect 530310 18359 530316 18367
rect 538142 18359 538148 18366
rect 530310 18323 538148 18359
rect 530310 18315 530316 18323
rect 538142 18314 538148 18323
rect 538200 18359 538206 18366
rect 538200 18323 538213 18359
rect 538200 18314 538206 18323
rect 530168 18275 530174 18283
rect 530166 18239 530174 18275
rect 530168 18231 530174 18239
rect 530226 18275 530232 18283
rect 538030 18275 538036 18282
rect 530226 18239 538036 18275
rect 530226 18231 530232 18239
rect 538030 18230 538036 18239
rect 538088 18275 538094 18282
rect 538088 18239 538101 18275
rect 538088 18230 538094 18239
rect 530084 18191 530090 18199
rect 530082 18155 530090 18191
rect 530084 18147 530090 18155
rect 530142 18191 530148 18199
rect 537918 18191 537924 18198
rect 530142 18155 537924 18191
rect 530142 18147 530148 18155
rect 537918 18146 537924 18155
rect 537976 18191 537982 18198
rect 537976 18155 537989 18191
rect 537976 18146 537982 18155
rect 530000 18107 530006 18115
rect 529998 18071 530006 18107
rect 530000 18063 530006 18071
rect 530058 18107 530064 18115
rect 537806 18107 537812 18114
rect 530058 18071 537812 18107
rect 530058 18063 530064 18071
rect 537806 18062 537812 18071
rect 537864 18107 537870 18114
rect 537864 18071 537877 18107
rect 537864 18062 537870 18071
rect 529916 18023 529922 18031
rect 529914 17987 529922 18023
rect 529916 17979 529922 17987
rect 529974 18023 529980 18031
rect 537694 18023 537700 18030
rect 529974 17987 537700 18023
rect 529974 17979 529980 17987
rect 537694 17978 537700 17987
rect 537752 18023 537758 18030
rect 537752 17987 537765 18023
rect 537752 17978 537758 17987
rect 529832 17939 529838 17947
rect 529830 17903 529838 17939
rect 529832 17895 529838 17903
rect 529890 17939 529896 17947
rect 537582 17939 537588 17946
rect 529890 17903 537588 17939
rect 529890 17895 529896 17903
rect 537582 17894 537588 17903
rect 537640 17939 537646 17946
rect 537640 17903 537653 17939
rect 537640 17894 537646 17903
rect 529748 17855 529754 17863
rect 529746 17819 529754 17855
rect 529748 17811 529754 17819
rect 529806 17855 529812 17863
rect 537470 17855 537476 17862
rect 529806 17819 537476 17855
rect 529806 17811 529812 17819
rect 537470 17810 537476 17819
rect 537528 17855 537534 17862
rect 537528 17819 537541 17855
rect 537528 17810 537534 17819
rect 529664 17771 529670 17779
rect 529662 17735 529670 17771
rect 529664 17727 529670 17735
rect 529722 17771 529728 17779
rect 537358 17771 537364 17778
rect 529722 17735 537364 17771
rect 529722 17727 529728 17735
rect 537358 17726 537364 17735
rect 537416 17771 537422 17778
rect 537416 17735 537429 17771
rect 537416 17726 537422 17735
rect 529580 17687 529586 17695
rect 529578 17651 529586 17687
rect 529580 17643 529586 17651
rect 529638 17687 529644 17695
rect 537246 17687 537252 17694
rect 529638 17651 537252 17687
rect 529638 17643 529644 17651
rect 537246 17642 537252 17651
rect 537304 17687 537310 17694
rect 537304 17651 537317 17687
rect 537304 17642 537310 17651
rect 529496 17603 529502 17611
rect 529494 17567 529502 17603
rect 529496 17559 529502 17567
rect 529554 17603 529560 17611
rect 537134 17603 537140 17610
rect 529554 17567 537140 17603
rect 529554 17559 529560 17567
rect 537134 17558 537140 17567
rect 537192 17603 537198 17610
rect 537192 17567 537205 17603
rect 537192 17558 537198 17567
rect 529412 17519 529418 17527
rect 529410 17483 529418 17519
rect 529412 17475 529418 17483
rect 529470 17519 529476 17527
rect 537022 17519 537028 17526
rect 529470 17483 537028 17519
rect 529470 17475 529476 17483
rect 537022 17474 537028 17483
rect 537080 17519 537086 17526
rect 537080 17483 537093 17519
rect 537080 17474 537086 17483
rect 529328 17435 529334 17443
rect 529326 17399 529334 17435
rect 529328 17391 529334 17399
rect 529386 17435 529392 17443
rect 536910 17435 536916 17442
rect 529386 17399 536916 17435
rect 529386 17391 529392 17399
rect 536910 17390 536916 17399
rect 536968 17435 536974 17442
rect 536968 17399 536981 17435
rect 536968 17390 536974 17399
rect 536686 17119 536692 17132
rect 520368 17083 536692 17119
rect 489074 9474 489110 11994
rect 490687 9798 490755 12012
rect 490687 9724 490755 9730
rect 520368 9474 520404 17083
rect 536686 17080 536692 17083
rect 536744 17080 536750 17132
rect 536574 17035 536580 17048
rect 520452 16999 536580 17035
rect 520452 11282 520488 16999
rect 536574 16996 536580 16999
rect 536632 16996 536638 17048
rect 536462 16951 536468 16964
rect 520536 16915 536468 16951
rect 520536 11402 520572 16915
rect 536462 16912 536468 16915
rect 536520 16912 536526 16964
rect 536350 16867 536356 16880
rect 520620 16831 536356 16867
rect 520620 11522 520656 16831
rect 536350 16828 536356 16831
rect 536408 16828 536414 16880
rect 536238 16783 536244 16796
rect 520704 16747 536244 16783
rect 520704 11642 520740 16747
rect 536238 16744 536244 16747
rect 536296 16744 536302 16796
rect 536126 16699 536132 16712
rect 520788 16663 536132 16699
rect 520788 13874 520824 16663
rect 536126 16660 536132 16663
rect 536184 16660 536190 16712
rect 536014 16615 536020 16628
rect 520872 16579 536020 16615
rect 520872 13994 520908 16579
rect 536014 16576 536020 16579
rect 536072 16576 536078 16628
rect 535902 16531 535908 16544
rect 520956 16495 535908 16531
rect 520956 14110 520992 16495
rect 535902 16492 535908 16495
rect 535960 16492 535966 16544
rect 535790 16447 535796 16460
rect 521040 16411 535796 16447
rect 521040 14234 521076 16411
rect 535790 16408 535796 16411
rect 535848 16408 535854 16460
rect 535678 16363 535684 16376
rect 521124 16327 535684 16363
rect 521032 14228 521084 14234
rect 521032 14170 521084 14176
rect 521040 14164 521076 14170
rect 520948 14104 521000 14110
rect 520948 14046 521000 14052
rect 520956 14042 520992 14046
rect 520860 13988 520912 13994
rect 520860 13930 520912 13936
rect 520872 13926 520908 13930
rect 520776 13868 520828 13874
rect 520776 13810 520828 13816
rect 520788 13804 520824 13810
rect 521124 13804 521160 16327
rect 535678 16324 535684 16327
rect 535736 16324 535742 16376
rect 535566 16279 535572 16292
rect 521208 16243 535572 16279
rect 521208 13804 521244 16243
rect 535566 16240 535572 16243
rect 535624 16240 535630 16292
rect 535454 16195 535460 16208
rect 521292 16159 535460 16195
rect 521292 13804 521328 16159
rect 535454 16156 535460 16159
rect 535512 16156 535518 16208
rect 535342 16111 535348 16124
rect 521376 16075 535348 16111
rect 521376 13804 521412 16075
rect 535342 16072 535348 16075
rect 535400 16072 535406 16124
rect 524412 15786 524418 15838
rect 524470 15830 524476 15838
rect 553374 15830 553380 15842
rect 524470 15794 553380 15830
rect 524470 15786 524476 15794
rect 553374 15790 553380 15794
rect 553432 15830 553438 15842
rect 553432 15794 553442 15830
rect 553432 15790 553438 15794
rect 524328 15702 524334 15754
rect 524386 15746 524392 15754
rect 553262 15746 553268 15756
rect 524386 15710 553268 15746
rect 524386 15702 524392 15710
rect 553262 15704 553268 15710
rect 553320 15746 553326 15756
rect 553320 15710 553334 15746
rect 553320 15704 553326 15710
rect 524244 15618 524250 15670
rect 524302 15662 524308 15670
rect 552926 15662 552932 15674
rect 524302 15626 552932 15662
rect 524302 15618 524308 15626
rect 552926 15622 552932 15626
rect 552984 15622 552990 15674
rect 524160 15534 524166 15586
rect 524218 15578 524224 15586
rect 552478 15578 552484 15592
rect 524218 15542 552484 15578
rect 524218 15534 524224 15542
rect 552478 15540 552484 15542
rect 552536 15578 552542 15592
rect 552536 15542 552544 15578
rect 552536 15540 552542 15542
rect 524076 15450 524082 15502
rect 524134 15494 524140 15502
rect 552142 15494 552148 15504
rect 524134 15458 552148 15494
rect 524134 15450 524140 15458
rect 552142 15452 552148 15458
rect 552200 15494 552206 15504
rect 552200 15458 552214 15494
rect 552200 15452 552206 15458
rect 523992 15366 523998 15418
rect 524050 15410 524056 15418
rect 551134 15410 551140 15422
rect 524050 15374 551140 15410
rect 524050 15366 524056 15374
rect 551134 15370 551140 15374
rect 551192 15410 551198 15422
rect 551192 15374 551200 15410
rect 551192 15370 551198 15374
rect 523908 15282 523914 15334
rect 523966 15326 523972 15334
rect 551022 15326 551028 15340
rect 523966 15290 551028 15326
rect 523966 15282 523972 15290
rect 551022 15288 551028 15290
rect 551080 15326 551086 15340
rect 551080 15290 551092 15326
rect 551080 15288 551086 15290
rect 523824 15198 523830 15250
rect 523882 15242 523888 15250
rect 550686 15242 550692 15254
rect 523882 15206 550692 15242
rect 523882 15198 523888 15206
rect 550686 15202 550692 15206
rect 550744 15242 550750 15254
rect 550744 15206 550754 15242
rect 550744 15202 550750 15206
rect 523740 15114 523746 15166
rect 523798 15158 523804 15166
rect 550126 15158 550132 15170
rect 523798 15122 550132 15158
rect 523798 15114 523804 15122
rect 550126 15118 550132 15122
rect 550184 15158 550190 15170
rect 550184 15122 550194 15158
rect 550184 15118 550190 15122
rect 523656 15030 523662 15082
rect 523714 15074 523720 15082
rect 549790 15074 549796 15092
rect 523714 15040 549796 15074
rect 549848 15074 549854 15092
rect 549848 15040 549856 15074
rect 523714 15038 549856 15040
rect 523714 15030 523720 15038
rect 523572 14946 523578 14998
rect 523630 14990 523636 14998
rect 545422 14990 545428 15006
rect 523630 14954 545428 14990
rect 545480 14990 545486 15006
rect 545480 14954 545490 14990
rect 523630 14946 523636 14954
rect 523488 14862 523494 14914
rect 523546 14906 523552 14914
rect 544638 14906 544644 14922
rect 523546 14870 544644 14906
rect 544696 14906 544702 14922
rect 544696 14870 544712 14906
rect 523546 14862 523552 14870
rect 523404 14778 523410 14830
rect 523462 14822 523468 14830
rect 543966 14822 543972 14832
rect 523462 14786 543972 14822
rect 523462 14778 523468 14786
rect 543966 14780 543972 14786
rect 544024 14822 544030 14832
rect 544024 14786 544034 14822
rect 544024 14780 544030 14786
rect 523320 14694 523326 14746
rect 523378 14738 523384 14746
rect 543182 14738 543188 14752
rect 523378 14702 543188 14738
rect 523378 14694 523384 14702
rect 543182 14700 543188 14702
rect 543240 14738 543246 14752
rect 543240 14702 543252 14738
rect 543240 14700 543246 14702
rect 529036 14436 529042 14444
rect 529023 14400 529042 14436
rect 529036 14392 529042 14400
rect 529094 14436 529100 14444
rect 529094 14400 555444 14436
rect 529094 14392 529100 14400
rect 528952 14362 528958 14370
rect 528939 14326 528958 14362
rect 528952 14318 528958 14326
rect 529010 14362 529016 14370
rect 529010 14326 555336 14362
rect 529010 14318 529016 14326
rect 528868 14288 528874 14296
rect 528855 14252 528874 14288
rect 528868 14244 528874 14252
rect 528926 14288 528932 14296
rect 528926 14252 555226 14288
rect 528926 14244 528932 14252
rect 528784 14214 528790 14222
rect 528771 14178 528790 14214
rect 528784 14170 528790 14178
rect 528842 14214 528848 14222
rect 528842 14178 554886 14214
rect 528842 14170 528848 14178
rect 528700 14140 528706 14148
rect 528687 14104 528706 14140
rect 528700 14096 528706 14104
rect 528758 14140 528764 14148
rect 528758 14104 554776 14140
rect 528758 14096 528764 14104
rect 528616 14066 528622 14074
rect 528603 14030 528622 14066
rect 528616 14022 528622 14030
rect 528674 14066 528680 14074
rect 528674 14030 553880 14066
rect 528674 14022 528680 14030
rect 528532 13992 528538 14000
rect 528519 13956 528538 13992
rect 528532 13948 528538 13956
rect 528590 13992 528596 14000
rect 528590 13956 553762 13992
rect 528590 13948 528596 13956
rect 528448 13918 528454 13926
rect 528435 13882 528454 13918
rect 528448 13874 528454 13882
rect 528506 13918 528512 13926
rect 528506 13882 553650 13918
rect 528506 13874 528512 13882
rect 528364 13844 528370 13852
rect 528351 13808 528370 13844
rect 528364 13800 528370 13808
rect 528422 13844 528428 13852
rect 528422 13808 552874 13844
rect 528422 13800 528428 13808
rect 528280 13770 528286 13778
rect 528267 13734 528286 13770
rect 528280 13726 528286 13734
rect 528338 13770 528344 13778
rect 528338 13734 552756 13770
rect 528338 13726 528344 13734
rect 528196 13696 528202 13704
rect 528183 13660 528202 13696
rect 528196 13652 528202 13660
rect 528254 13696 528260 13704
rect 528254 13660 551648 13696
rect 528254 13652 528260 13660
rect 528112 13622 528118 13630
rect 528099 13586 528118 13622
rect 528112 13578 528118 13586
rect 528170 13622 528176 13630
rect 528170 13586 551534 13622
rect 528170 13578 528176 13586
rect 528028 13548 528034 13556
rect 528015 13512 528034 13548
rect 528028 13504 528034 13512
rect 528086 13548 528092 13556
rect 528086 13512 551422 13548
rect 528086 13504 528092 13512
rect 527944 13474 527950 13482
rect 527931 13438 527950 13474
rect 527944 13430 527950 13438
rect 528002 13474 528008 13482
rect 528002 13438 550644 13474
rect 528002 13430 528008 13438
rect 527860 13400 527866 13408
rect 527847 13364 527866 13400
rect 527860 13356 527866 13364
rect 527918 13400 527924 13408
rect 527918 13364 550520 13400
rect 527918 13356 527924 13364
rect 527776 13326 527782 13334
rect 527763 13290 527782 13326
rect 527776 13282 527782 13290
rect 527834 13326 527840 13334
rect 527834 13290 550400 13326
rect 527834 13282 527840 13290
rect 527692 13252 527698 13260
rect 527679 13216 527698 13252
rect 527692 13208 527698 13216
rect 527750 13252 527756 13260
rect 527750 13216 549292 13252
rect 527750 13208 527756 13216
rect 527608 13178 527614 13186
rect 527595 13142 527614 13178
rect 527608 13134 527614 13142
rect 527666 13178 527672 13186
rect 527666 13142 549170 13178
rect 527666 13134 527672 13142
rect 527524 13104 527530 13112
rect 527511 13068 527530 13104
rect 527524 13060 527530 13068
rect 527582 13104 527588 13112
rect 527582 13068 549066 13104
rect 527582 13060 527588 13068
rect 527440 13030 527446 13038
rect 527427 12994 527446 13030
rect 527440 12986 527446 12994
rect 527498 13030 527504 13038
rect 527498 12994 548954 13030
rect 527498 12986 527504 12994
rect 527356 12956 527362 12964
rect 527343 12920 527362 12956
rect 527356 12912 527362 12920
rect 527414 12956 527420 12964
rect 527414 12920 548844 12956
rect 527414 12912 527420 12920
rect 527272 12882 527278 12890
rect 527259 12846 527278 12882
rect 527272 12838 527278 12846
rect 527330 12882 527336 12890
rect 527330 12846 548734 12882
rect 527330 12838 527336 12846
rect 527188 12808 527194 12816
rect 527175 12772 527194 12808
rect 527188 12764 527194 12772
rect 527246 12808 527252 12816
rect 527246 12772 548626 12808
rect 527246 12764 527252 12772
rect 527104 12734 527110 12742
rect 527091 12698 527110 12734
rect 527104 12690 527110 12698
rect 527162 12734 527168 12742
rect 527162 12698 548506 12734
rect 527162 12690 527168 12698
rect 527020 12660 527026 12668
rect 527007 12624 527026 12660
rect 527020 12616 527026 12624
rect 527078 12660 527084 12668
rect 527078 12624 548388 12660
rect 527078 12616 527084 12624
rect 526936 12586 526942 12594
rect 526923 12550 526942 12586
rect 526936 12542 526942 12550
rect 526994 12586 527000 12594
rect 526994 12550 548280 12586
rect 526994 12542 527000 12550
rect 526852 12512 526858 12520
rect 526839 12476 526858 12512
rect 526852 12468 526858 12476
rect 526910 12512 526916 12520
rect 526910 12476 548052 12512
rect 526910 12468 526916 12476
rect 526768 12438 526774 12446
rect 526755 12402 526774 12438
rect 526768 12394 526774 12402
rect 526826 12438 526832 12446
rect 526826 12402 547930 12438
rect 526826 12394 526832 12402
rect 526684 12364 526690 12372
rect 526671 12328 526690 12364
rect 526684 12320 526690 12328
rect 526742 12364 526748 12372
rect 526742 12328 547826 12364
rect 526742 12320 526748 12328
rect 526600 12290 526606 12298
rect 526587 12254 526606 12290
rect 526600 12246 526606 12254
rect 526658 12290 526664 12298
rect 526658 12254 547610 12290
rect 526658 12246 526664 12254
rect 526516 12216 526522 12224
rect 526503 12180 526522 12216
rect 526516 12172 526522 12180
rect 526574 12216 526580 12224
rect 526574 12180 547502 12216
rect 526574 12172 526580 12180
rect 526432 12142 526438 12150
rect 526419 12106 526438 12142
rect 526432 12098 526438 12106
rect 526490 12142 526496 12150
rect 526490 12106 547274 12142
rect 526490 12098 526496 12106
rect 526348 12068 526354 12076
rect 526335 12032 526354 12068
rect 526348 12024 526354 12032
rect 526406 12068 526412 12076
rect 526406 12032 547164 12068
rect 526406 12024 526412 12032
rect 526264 11994 526270 12002
rect 526251 11958 526270 11994
rect 526264 11950 526270 11958
rect 526322 11994 526328 12002
rect 526322 11958 547048 11994
rect 526322 11950 526328 11958
rect 526180 11920 526186 11928
rect 526167 11884 526186 11920
rect 526180 11876 526186 11884
rect 526238 11920 526244 11928
rect 526238 11884 546824 11920
rect 526238 11876 526244 11884
rect 526096 11846 526102 11854
rect 526083 11810 526102 11846
rect 526096 11802 526102 11810
rect 526154 11846 526160 11854
rect 526154 11810 546722 11846
rect 526154 11802 526160 11810
rect 526012 11772 526018 11780
rect 525999 11736 526018 11772
rect 526012 11728 526018 11736
rect 526070 11772 526076 11780
rect 526070 11736 546594 11772
rect 526070 11728 526076 11736
rect 525928 11698 525934 11706
rect 525915 11662 525934 11698
rect 525928 11654 525934 11662
rect 525986 11698 525992 11706
rect 525986 11662 546384 11698
rect 525986 11654 525992 11662
rect 520698 11636 520750 11642
rect 525844 11624 525850 11632
rect 525831 11588 525850 11624
rect 520698 11578 520750 11584
rect 525844 11580 525850 11588
rect 525902 11624 525908 11632
rect 525902 11588 546256 11624
rect 525902 11580 525908 11588
rect 520704 11572 520740 11578
rect 525760 11550 525766 11558
rect 520612 11516 520664 11522
rect 525747 11514 525766 11550
rect 525760 11506 525766 11514
rect 525818 11550 525824 11558
rect 525818 11514 546042 11550
rect 525818 11506 525824 11514
rect 525676 11476 525682 11484
rect 520612 11458 520664 11464
rect 520620 11454 520656 11458
rect 525663 11440 525682 11476
rect 525676 11432 525682 11440
rect 525734 11476 525740 11484
rect 525734 11440 545926 11476
rect 525734 11432 525740 11440
rect 525592 11402 525598 11410
rect 520526 11396 520578 11402
rect 525579 11366 525598 11402
rect 525592 11358 525598 11366
rect 525650 11402 525656 11410
rect 525650 11366 545816 11402
rect 525650 11358 525656 11366
rect 520526 11338 520578 11344
rect 525508 11328 525514 11336
rect 525495 11292 525514 11328
rect 525508 11284 525514 11292
rect 525566 11328 525572 11336
rect 525566 11292 545378 11328
rect 525566 11284 525572 11292
rect 520442 11276 520494 11282
rect 525424 11254 525430 11262
rect 520442 11218 520494 11224
rect 525411 11218 525430 11254
rect 520452 11210 520488 11218
rect 525424 11210 525430 11218
rect 525482 11254 525488 11262
rect 525482 11218 545254 11254
rect 525482 11210 525488 11218
rect 525340 11180 525346 11188
rect 525327 11144 525346 11180
rect 525340 11136 525346 11144
rect 525398 11180 525404 11188
rect 525398 11144 545140 11180
rect 525398 11136 525404 11144
rect 525256 11106 525262 11114
rect 525243 11070 525262 11106
rect 525256 11062 525262 11070
rect 525314 11106 525320 11114
rect 525314 11070 545030 11106
rect 525314 11062 525320 11070
rect 525172 11032 525178 11040
rect 525159 10996 525178 11032
rect 525172 10988 525178 10996
rect 525230 11032 525236 11040
rect 525230 10996 544588 11032
rect 525230 10988 525236 10996
rect 525088 10958 525094 10966
rect 525075 10922 525094 10958
rect 525088 10914 525094 10922
rect 525146 10958 525152 10966
rect 525146 10922 544476 10958
rect 525146 10914 525152 10922
rect 525004 10884 525010 10892
rect 524991 10848 525010 10884
rect 525004 10840 525010 10848
rect 525062 10884 525068 10892
rect 525062 10848 544352 10884
rect 525062 10840 525068 10848
rect 524920 10810 524926 10818
rect 524907 10774 524926 10810
rect 524920 10766 524926 10774
rect 524978 10810 524984 10818
rect 524978 10774 543920 10810
rect 524978 10766 524984 10774
rect 524836 10736 524842 10744
rect 524823 10700 524842 10736
rect 524836 10692 524842 10700
rect 524894 10736 524900 10744
rect 524894 10700 543808 10736
rect 524894 10692 524900 10700
rect 524752 10662 524758 10670
rect 524739 10626 524758 10662
rect 524752 10618 524758 10626
rect 524810 10662 524816 10670
rect 524810 10626 543692 10662
rect 524810 10618 524816 10626
rect 524668 10588 524674 10596
rect 524655 10552 524674 10588
rect 524668 10544 524674 10552
rect 524726 10588 524732 10596
rect 524726 10552 543576 10588
rect 524726 10544 524732 10552
rect 534782 10367 534788 10380
rect 489074 9438 520404 9474
rect 521611 10331 534788 10367
rect 521611 9369 521647 10331
rect 534782 10328 534788 10331
rect 534840 10367 534846 10380
rect 534840 10331 534855 10367
rect 534840 10328 534846 10331
rect 535236 10295 535288 10301
rect 483820 9333 521647 9369
rect 521695 10247 535236 10283
rect 521695 9285 521731 10247
rect 535288 10247 535301 10283
rect 535236 10237 535288 10243
rect 535118 10199 535124 10211
rect 483736 9249 521731 9285
rect 521779 10163 535124 10199
rect 521779 9201 521815 10163
rect 535118 10159 535124 10163
rect 535176 10199 535182 10211
rect 535176 10163 535191 10199
rect 535176 10159 535182 10163
rect 535006 10115 535012 10127
rect 483652 9165 521815 9201
rect 521863 10079 535012 10115
rect 521863 9117 521899 10079
rect 535006 10075 535012 10079
rect 535064 10115 535070 10127
rect 535064 10079 535084 10115
rect 535064 10075 535070 10079
rect 534894 10031 534900 10041
rect 483568 9081 521899 9117
rect 521947 9995 534900 10031
rect 521947 9033 521983 9995
rect 534894 9989 534900 9995
rect 534952 10031 534958 10041
rect 534952 9995 534966 10031
rect 534952 9989 534958 9995
rect 522949 9921 522955 9930
rect 522945 9885 522955 9921
rect 522949 9878 522955 9885
rect 523007 9921 523013 9930
rect 539934 9921 539940 9932
rect 523007 9885 539940 9921
rect 523007 9878 523013 9885
rect 539934 9880 539940 9885
rect 539992 9921 539998 9932
rect 539992 9885 540012 9921
rect 539992 9880 539998 9885
rect 522865 9837 522871 9846
rect 522861 9801 522871 9837
rect 522865 9794 522871 9801
rect 522923 9837 522929 9846
rect 539822 9837 539828 9848
rect 522923 9801 539828 9837
rect 522923 9794 522929 9801
rect 539822 9796 539828 9801
rect 539880 9837 539886 9848
rect 539880 9801 539900 9837
rect 539880 9796 539886 9801
rect 522781 9753 522787 9762
rect 522777 9717 522787 9753
rect 522781 9710 522787 9717
rect 522839 9753 522845 9762
rect 539710 9753 539716 9764
rect 522839 9717 539716 9753
rect 522839 9710 522845 9717
rect 539710 9712 539716 9717
rect 539768 9753 539774 9764
rect 539768 9717 539788 9753
rect 539768 9712 539774 9717
rect 522697 9669 522703 9678
rect 522693 9633 522703 9669
rect 522697 9626 522703 9633
rect 522755 9669 522761 9678
rect 539598 9669 539604 9680
rect 522755 9633 539604 9669
rect 522755 9626 522761 9633
rect 539598 9628 539604 9633
rect 539656 9669 539662 9680
rect 539656 9633 539676 9669
rect 539656 9628 539662 9633
rect 522613 9585 522619 9594
rect 522609 9549 522619 9585
rect 522613 9542 522619 9549
rect 522671 9585 522677 9594
rect 539486 9585 539492 9596
rect 522671 9549 539492 9585
rect 522671 9542 522677 9549
rect 539486 9544 539492 9549
rect 539544 9585 539550 9596
rect 539544 9549 539564 9585
rect 539544 9544 539550 9549
rect 522529 9501 522535 9510
rect 522525 9465 522535 9501
rect 522529 9458 522535 9465
rect 522587 9501 522593 9510
rect 539374 9501 539380 9512
rect 522587 9465 539380 9501
rect 522587 9458 522593 9465
rect 539374 9460 539380 9465
rect 539432 9501 539438 9512
rect 539432 9465 539452 9501
rect 539432 9460 539438 9465
rect 522445 9417 522451 9426
rect 522441 9381 522451 9417
rect 522445 9374 522451 9381
rect 522503 9417 522509 9426
rect 539262 9417 539268 9428
rect 522503 9381 539268 9417
rect 522503 9374 522509 9381
rect 539262 9376 539268 9381
rect 539320 9417 539326 9428
rect 539320 9381 539340 9417
rect 539320 9376 539326 9381
rect 522361 9333 522367 9342
rect 522357 9297 522367 9333
rect 522361 9290 522367 9297
rect 522419 9333 522425 9342
rect 539150 9333 539156 9344
rect 522419 9297 539156 9333
rect 522419 9290 522425 9297
rect 539150 9292 539156 9297
rect 539208 9333 539214 9344
rect 539208 9297 539228 9333
rect 539208 9292 539214 9297
rect 522277 9249 522283 9258
rect 522273 9213 522283 9249
rect 522277 9206 522283 9213
rect 522335 9249 522341 9258
rect 539038 9249 539044 9260
rect 522335 9213 539044 9249
rect 522335 9206 522341 9213
rect 539038 9208 539044 9213
rect 539096 9249 539102 9260
rect 539096 9213 539116 9249
rect 539096 9208 539102 9213
rect 522193 9165 522199 9174
rect 522189 9129 522199 9165
rect 522193 9122 522199 9129
rect 522251 9165 522257 9174
rect 538926 9165 538932 9176
rect 522251 9129 538932 9165
rect 522251 9122 522257 9129
rect 538926 9124 538932 9129
rect 538984 9165 538990 9176
rect 538984 9129 539004 9165
rect 538984 9124 538990 9129
rect 522109 9081 522115 9090
rect 522105 9045 522115 9081
rect 522109 9038 522115 9045
rect 522167 9081 522173 9090
rect 538814 9081 538820 9092
rect 522167 9045 538820 9081
rect 522167 9038 522173 9045
rect 538814 9040 538820 9045
rect 538872 9081 538878 9092
rect 538872 9045 538892 9081
rect 538872 9040 538878 9045
rect 25374 9018 25380 9031
rect 25372 8982 25380 9018
rect 25374 8979 25380 8982
rect 25432 9018 25438 9031
rect 98344 9018 98350 9023
rect 25432 8982 98350 9018
rect 25432 8979 25438 8982
rect 98344 8971 98350 8982
rect 98402 9018 98408 9023
rect 98402 8982 98416 9018
rect 483484 8997 521983 9033
rect 522025 8997 522031 9006
rect 98402 8971 98408 8982
rect 522021 8961 522031 8997
rect 522025 8954 522031 8961
rect 522083 8997 522089 9006
rect 538702 8997 538708 9008
rect 522083 8961 538708 8997
rect 522083 8954 522089 8961
rect 538702 8956 538708 8961
rect 538760 8997 538766 9008
rect 538760 8961 538780 8997
rect 538760 8956 538766 8961
rect 25492 8947 25544 8953
rect 25484 8898 25492 8934
rect 99972 8934 99978 8939
rect 25544 8898 99978 8934
rect 25492 8889 25544 8895
rect 99972 8887 99978 8898
rect 100030 8934 100036 8939
rect 100030 8898 100043 8934
rect 521941 8913 521947 8922
rect 100030 8887 100036 8898
rect 521937 8877 521947 8913
rect 521941 8870 521947 8877
rect 521999 8913 522005 8922
rect 538590 8913 538596 8924
rect 521999 8877 538596 8913
rect 521999 8870 522005 8877
rect 538590 8872 538596 8877
rect 538648 8913 538654 8924
rect 538648 8877 538668 8913
rect 538648 8872 538654 8877
rect 25598 8850 25604 8863
rect 25596 8814 25604 8850
rect 25598 8811 25604 8814
rect 25656 8850 25662 8863
rect 101600 8850 101606 8855
rect 25656 8814 101606 8850
rect 25656 8811 25662 8814
rect 101600 8803 101606 8814
rect 101658 8850 101664 8855
rect 101658 8814 101672 8850
rect 521857 8829 521863 8838
rect 101658 8803 101664 8814
rect 521853 8793 521863 8829
rect 521857 8786 521863 8793
rect 521915 8829 521921 8838
rect 538478 8829 538484 8840
rect 521915 8793 538484 8829
rect 521915 8786 521921 8793
rect 538478 8788 538484 8793
rect 538536 8829 538542 8840
rect 538536 8793 538556 8829
rect 538536 8788 538542 8793
rect 25710 8766 25716 8779
rect 25708 8730 25716 8766
rect 25710 8727 25716 8730
rect 25768 8766 25774 8779
rect 103228 8766 103234 8771
rect 25768 8730 103234 8766
rect 25768 8727 25774 8730
rect 103228 8719 103234 8730
rect 103286 8766 103292 8771
rect 103286 8730 103296 8766
rect 521773 8745 521779 8754
rect 103286 8719 103292 8730
rect 521769 8709 521779 8745
rect 521773 8702 521779 8709
rect 521831 8745 521837 8754
rect 538366 8745 538372 8756
rect 521831 8709 538372 8745
rect 521831 8702 521837 8709
rect 538366 8704 538372 8709
rect 538424 8745 538430 8756
rect 538424 8709 538444 8745
rect 538424 8704 538430 8709
rect 25822 8682 25828 8696
rect 25820 8646 25828 8682
rect 25822 8644 25828 8646
rect 25880 8682 25886 8696
rect 104856 8682 104862 8693
rect 25880 8646 104862 8682
rect 25880 8644 25886 8646
rect 104856 8641 104862 8646
rect 104914 8682 104920 8693
rect 104914 8646 104923 8682
rect 521689 8661 521695 8670
rect 104914 8641 104920 8646
rect 521685 8625 521695 8661
rect 521689 8618 521695 8625
rect 521747 8661 521753 8670
rect 538254 8661 538260 8671
rect 521747 8625 538260 8661
rect 521747 8618 521753 8625
rect 538254 8619 538260 8625
rect 538312 8661 538318 8671
rect 538312 8625 538332 8661
rect 538312 8619 538318 8625
rect 484686 8524 484692 8532
rect 484676 8488 484692 8524
rect 484686 8480 484692 8488
rect 484744 8524 484750 8532
rect 542616 8524 542622 8532
rect 484744 8488 542622 8524
rect 484744 8480 484750 8488
rect 542616 8480 542622 8488
rect 542674 8480 542680 8532
rect 484602 8440 484608 8448
rect 484592 8404 484608 8440
rect 484602 8396 484608 8404
rect 484660 8440 484666 8448
rect 542504 8440 542510 8448
rect 484660 8404 542510 8440
rect 484660 8396 484666 8404
rect 542504 8396 542510 8404
rect 542562 8440 542568 8448
rect 542562 8404 542576 8440
rect 542562 8396 542568 8404
rect 484518 8356 484524 8364
rect 484508 8320 484524 8356
rect 484518 8312 484524 8320
rect 484576 8356 484582 8364
rect 542392 8356 542398 8364
rect 484576 8320 542398 8356
rect 484576 8312 484582 8320
rect 542392 8312 542398 8320
rect 542450 8312 542458 8364
rect 484434 8272 484440 8280
rect 484424 8236 484440 8272
rect 484434 8228 484440 8236
rect 484492 8272 484498 8280
rect 542280 8272 542286 8280
rect 484492 8236 542286 8272
rect 484492 8228 484498 8236
rect 542280 8228 542286 8236
rect 542338 8272 542344 8280
rect 542338 8236 542346 8272
rect 542338 8228 542344 8236
rect 484350 8188 484356 8196
rect 484340 8152 484356 8188
rect 484350 8144 484356 8152
rect 484408 8188 484414 8196
rect 542168 8188 542174 8196
rect 484408 8152 542174 8188
rect 484408 8144 484414 8152
rect 542168 8144 542174 8152
rect 542226 8188 542232 8196
rect 542226 8152 542236 8188
rect 542226 8144 542232 8152
rect 484266 8104 484272 8112
rect 484256 8068 484272 8104
rect 484266 8060 484272 8068
rect 484324 8104 484330 8112
rect 542056 8104 542062 8112
rect 484324 8068 542062 8104
rect 484324 8060 484330 8068
rect 542056 8060 542062 8068
rect 542114 8104 542120 8112
rect 542114 8068 542126 8104
rect 542114 8060 542120 8068
rect 484182 8020 484188 8028
rect 484172 7984 484188 8020
rect 484182 7976 484188 7984
rect 484240 8020 484246 8028
rect 541944 8020 541950 8028
rect 484240 7984 541950 8020
rect 484240 7976 484246 7984
rect 541944 7976 541950 7984
rect 542002 8020 542008 8028
rect 542002 7984 542014 8020
rect 542002 7976 542008 7984
rect 484098 7936 484104 7944
rect 484088 7900 484104 7936
rect 484098 7892 484104 7900
rect 484156 7936 484162 7944
rect 541832 7936 541838 7944
rect 484156 7900 541838 7936
rect 484156 7892 484162 7900
rect 541832 7892 541838 7900
rect 541890 7936 541896 7944
rect 541890 7900 541910 7936
rect 541890 7892 541896 7900
rect 25934 7858 25940 7872
rect 25932 7822 25940 7858
rect 25934 7820 25940 7822
rect 25992 7858 25998 7872
rect 233036 7858 233042 7866
rect 25992 7822 233042 7858
rect 25992 7820 25998 7822
rect 233036 7814 233042 7822
rect 233094 7814 233100 7866
rect 484014 7852 484020 7860
rect 484004 7816 484020 7852
rect 484014 7808 484020 7816
rect 484072 7852 484078 7860
rect 541720 7852 541726 7860
rect 484072 7816 541726 7852
rect 484072 7808 484078 7816
rect 541720 7808 541726 7816
rect 541778 7852 541784 7860
rect 541778 7816 541790 7852
rect 541778 7808 541784 7816
rect 26046 7774 26052 7788
rect 26044 7738 26052 7774
rect 26046 7736 26052 7738
rect 26104 7774 26110 7788
rect 173946 7774 173952 7782
rect 26104 7738 173952 7774
rect 26104 7736 26110 7738
rect 173946 7730 173952 7738
rect 174004 7730 174010 7782
rect 483930 7768 483936 7776
rect 483920 7732 483936 7768
rect 483930 7724 483936 7732
rect 483988 7768 483994 7776
rect 541612 7768 541618 7776
rect 483988 7732 541618 7768
rect 483988 7724 483994 7732
rect 541612 7724 541618 7732
rect 541670 7724 541676 7776
rect 483846 7684 483852 7692
rect 483836 7648 483852 7684
rect 483846 7640 483852 7648
rect 483904 7684 483910 7692
rect 541504 7684 541510 7692
rect 483904 7648 541510 7684
rect 483904 7640 483910 7648
rect 541504 7640 541510 7648
rect 541562 7684 541568 7692
rect 541562 7648 541570 7684
rect 541562 7640 541568 7648
rect 483762 7600 483768 7608
rect 483752 7564 483768 7600
rect 483762 7556 483768 7564
rect 483820 7600 483826 7608
rect 541396 7600 541402 7608
rect 483820 7564 541402 7600
rect 483820 7556 483826 7564
rect 541396 7556 541402 7564
rect 541454 7600 541460 7608
rect 541454 7564 541472 7600
rect 541454 7556 541460 7564
rect 483678 7516 483684 7524
rect 483668 7480 483684 7516
rect 483678 7472 483684 7480
rect 483736 7516 483742 7524
rect 541284 7516 541290 7524
rect 483736 7480 541290 7516
rect 483736 7472 483742 7480
rect 541284 7472 541290 7480
rect 541342 7516 541348 7524
rect 541342 7480 541358 7516
rect 541342 7472 541348 7480
rect 483594 7432 483600 7440
rect 483584 7396 483600 7432
rect 483594 7388 483600 7396
rect 483652 7432 483658 7440
rect 541172 7432 541178 7440
rect 483652 7396 541178 7432
rect 483652 7388 483658 7396
rect 541172 7388 541178 7396
rect 541230 7432 541236 7440
rect 541230 7396 541246 7432
rect 541230 7388 541236 7396
rect 483510 7348 483516 7356
rect 483496 7312 483516 7348
rect 483510 7304 483516 7312
rect 483568 7348 483574 7356
rect 541060 7348 541066 7356
rect 483568 7312 541066 7348
rect 483568 7304 483574 7312
rect 541060 7304 541066 7312
rect 541118 7348 541124 7356
rect 541118 7312 541130 7348
rect 541118 7304 541124 7312
rect 483426 7264 483432 7272
rect 483420 7228 483432 7264
rect 483426 7220 483432 7228
rect 483484 7264 483490 7272
rect 540948 7264 540954 7272
rect 483484 7228 540954 7264
rect 483484 7220 483490 7228
rect 540948 7220 540954 7228
rect 541006 7264 541012 7272
rect 541006 7228 541022 7264
rect 541006 7220 541012 7228
rect 483342 7180 483348 7188
rect 483338 7144 483348 7180
rect 483342 7136 483348 7144
rect 483400 7180 483406 7188
rect 540834 7180 540840 7188
rect 483400 7144 540840 7180
rect 483400 7136 483406 7144
rect 540834 7136 540840 7144
rect 540892 7180 540898 7188
rect 540892 7144 540906 7180
rect 540892 7136 540898 7144
rect 483258 7096 483264 7104
rect 483248 7060 483264 7096
rect 483258 7052 483264 7060
rect 483316 7096 483322 7104
rect 540720 7096 540726 7104
rect 483316 7060 540726 7096
rect 483316 7052 483322 7060
rect 540720 7052 540726 7060
rect 540778 7052 540784 7104
rect 483174 7012 483180 7020
rect 483168 6976 483180 7012
rect 483174 6968 483180 6976
rect 483232 7012 483238 7020
rect 540606 7012 540612 7020
rect 483232 6976 540612 7012
rect 483232 6968 483238 6976
rect 540606 6968 540612 6976
rect 540664 7012 540670 7020
rect 540664 6976 540680 7012
rect 540664 6968 540670 6976
rect 483090 6928 483096 6936
rect 483086 6892 483096 6928
rect 483090 6884 483096 6892
rect 483148 6928 483154 6936
rect 540492 6928 540498 6936
rect 483148 6892 540498 6928
rect 483148 6884 483154 6892
rect 540492 6884 540498 6892
rect 540550 6928 540556 6936
rect 540550 6892 540564 6928
rect 540550 6884 540556 6892
rect 483006 6800 483012 6852
rect 483064 6844 483070 6852
rect 540378 6844 540384 6852
rect 483064 6808 540384 6844
rect 483064 6800 483070 6808
rect 540378 6800 540384 6808
rect 540436 6844 540442 6852
rect 540436 6808 540456 6844
rect 540436 6800 540442 6808
rect 17310 6726 17316 6778
rect 17368 6769 17374 6778
rect 34590 6769 34596 6778
rect 17368 6733 34596 6769
rect 17368 6726 17374 6733
rect 34590 6726 34596 6733
rect 34648 6769 34654 6778
rect 34648 6733 34657 6769
rect 34648 6726 34654 6733
rect 17646 6685 17652 6693
rect 17636 6649 17652 6685
rect 17646 6641 17652 6649
rect 17704 6685 17710 6693
rect 34674 6685 34680 6694
rect 17704 6649 34680 6685
rect 17704 6641 17710 6649
rect 34674 6642 34680 6649
rect 34732 6685 34738 6694
rect 34732 6649 34741 6685
rect 34732 6642 34738 6649
rect 17758 6601 17764 6608
rect 17745 6565 17764 6601
rect 17758 6556 17764 6565
rect 17816 6601 17822 6608
rect 34758 6601 34764 6610
rect 17816 6565 34764 6601
rect 17816 6556 17822 6565
rect 34758 6558 34764 6565
rect 34816 6601 34822 6610
rect 34816 6565 34825 6601
rect 34816 6558 34822 6565
rect 18094 6517 18100 6524
rect 18086 6481 18100 6517
rect 18094 6472 18100 6481
rect 18152 6517 18158 6524
rect 34842 6517 34848 6526
rect 18152 6481 34848 6517
rect 18152 6472 18158 6481
rect 34842 6474 34848 6481
rect 34900 6517 34906 6526
rect 34900 6481 34909 6517
rect 34900 6474 34906 6481
rect 18206 6433 18212 6440
rect 18196 6397 18212 6433
rect 18206 6388 18212 6397
rect 18264 6433 18270 6440
rect 34926 6433 34932 6442
rect 18264 6397 34932 6433
rect 18264 6388 18270 6397
rect 34926 6390 34932 6397
rect 34984 6433 34990 6442
rect 34984 6397 34993 6433
rect 34984 6390 34990 6397
rect 19438 6349 19444 6356
rect 19426 6313 19444 6349
rect 19438 6304 19444 6313
rect 19496 6349 19502 6356
rect 35010 6349 35016 6358
rect 19496 6313 35016 6349
rect 19496 6304 19502 6313
rect 35010 6306 35016 6313
rect 35068 6349 35074 6358
rect 35068 6313 35077 6349
rect 35068 6306 35074 6313
rect 19774 6265 19780 6274
rect 19762 6229 19780 6265
rect 19774 6222 19780 6229
rect 19832 6265 19838 6274
rect 35094 6265 35100 6274
rect 19832 6229 35100 6265
rect 19832 6222 19838 6229
rect 35094 6222 35100 6229
rect 35152 6265 35158 6274
rect 35152 6229 35161 6265
rect 35152 6222 35158 6229
rect 19886 6181 19892 6185
rect 19869 6145 19892 6181
rect 19886 6133 19892 6145
rect 19944 6181 19950 6185
rect 35178 6181 35184 6190
rect 19944 6145 35184 6181
rect 19944 6133 19950 6145
rect 35178 6138 35184 6145
rect 35236 6181 35242 6190
rect 35236 6145 35245 6181
rect 35236 6138 35242 6145
rect 20222 6097 20228 6102
rect 20216 6061 20228 6097
rect 20222 6050 20228 6061
rect 20280 6097 20286 6102
rect 35262 6097 35268 6106
rect 20280 6061 35268 6097
rect 20280 6050 20286 6061
rect 35262 6054 35268 6061
rect 35320 6097 35326 6106
rect 35320 6061 35329 6097
rect 35320 6054 35326 6061
rect 20334 6013 20340 6022
rect 20323 5977 20340 6013
rect 20334 5970 20340 5977
rect 20392 6013 20398 6022
rect 35346 6013 35352 6022
rect 20392 5977 35352 6013
rect 20392 5970 20398 5977
rect 35346 5970 35352 5977
rect 35404 6013 35410 6022
rect 35404 5977 35413 6013
rect 35404 5970 35410 5977
rect 20894 5929 20900 5939
rect 20883 5893 20900 5929
rect 20894 5887 20900 5893
rect 20952 5929 20958 5939
rect 35430 5929 35436 5938
rect 20952 5893 35436 5929
rect 20952 5887 20958 5893
rect 35430 5886 35436 5893
rect 35488 5929 35494 5938
rect 35488 5893 35497 5929
rect 35488 5886 35494 5893
rect 21118 5845 21124 5854
rect 21103 5809 21124 5845
rect 21118 5802 21124 5809
rect 21176 5845 21182 5854
rect 35514 5845 35520 5854
rect 21176 5809 35520 5845
rect 21176 5802 21182 5809
rect 35514 5802 35520 5809
rect 35572 5845 35578 5854
rect 35572 5809 35581 5845
rect 35572 5802 35578 5809
rect 13278 5565 13284 5617
rect 13336 5604 13342 5617
rect 13336 5568 94721 5604
rect 13336 5565 13342 5568
rect 13390 5480 13396 5532
rect 13448 5520 13454 5532
rect 13448 5484 94637 5520
rect 13448 5480 13454 5484
rect 13502 5396 13508 5448
rect 13560 5436 13566 5448
rect 13560 5400 94553 5436
rect 13560 5396 13566 5400
rect 13614 5312 13620 5364
rect 13672 5352 13678 5364
rect 13672 5316 94469 5352
rect 13672 5312 13678 5316
rect 13726 5268 13732 5280
rect 13725 5232 13732 5268
rect 13726 5228 13732 5232
rect 13784 5268 13790 5280
rect 13784 5232 94385 5268
rect 13784 5228 13790 5232
rect 13838 5145 13844 5197
rect 13896 5184 13902 5197
rect 13896 5148 94301 5184
rect 13896 5145 13902 5148
rect 15966 5060 15972 5112
rect 16024 5100 16030 5112
rect 16024 5064 94217 5100
rect 16024 5060 16030 5064
rect 16078 4978 16084 5030
rect 16136 5016 16142 5030
rect 16136 4980 94133 5016
rect 16136 4978 16142 4980
rect 16862 4932 16868 4946
rect 16858 4896 16868 4932
rect 16862 4894 16868 4896
rect 16920 4932 16926 4946
rect 16920 4896 94049 4932
rect 16920 4894 16926 4896
rect 16974 4808 16980 4860
rect 17032 4848 17038 4860
rect 17032 4812 93965 4848
rect 17032 4808 17038 4812
rect 17086 4723 17092 4775
rect 17144 4764 17150 4775
rect 17144 4728 93881 4764
rect 17144 4723 17150 4728
rect 17198 4642 17204 4694
rect 17256 4680 17262 4694
rect 17256 4644 93797 4680
rect 17256 4642 17262 4644
rect 17422 4557 17428 4609
rect 17480 4596 17486 4609
rect 17480 4560 93713 4596
rect 17480 4557 17486 4560
rect 17534 4473 17540 4525
rect 17592 4512 17598 4525
rect 17592 4476 93629 4512
rect 17592 4473 17598 4476
rect 17870 4305 17876 4357
rect 17928 4344 17934 4357
rect 17928 4308 93461 4344
rect 17928 4305 17934 4308
rect 17982 4220 17988 4272
rect 18040 4260 18046 4272
rect 18040 4224 93377 4260
rect 18040 4220 18046 4224
rect 18990 4136 18996 4188
rect 19048 4176 19054 4188
rect 19048 4140 93293 4176
rect 19048 4136 19054 4140
rect 19102 4053 19108 4105
rect 19160 4092 19166 4105
rect 19160 4056 93209 4092
rect 19160 4053 19166 4056
rect 19214 4008 19220 4021
rect 19212 3972 19220 4008
rect 19214 3969 19220 3972
rect 19272 4008 19278 4021
rect 19272 3972 93125 4008
rect 19272 3969 19278 3972
rect 19326 3885 19332 3937
rect 19384 3924 19390 3937
rect 19384 3888 93041 3924
rect 19384 3885 19390 3888
rect 19550 3840 19556 3854
rect 19544 3804 19556 3840
rect 19550 3802 19556 3804
rect 19608 3840 19614 3854
rect 19608 3804 92957 3840
rect 19608 3802 19614 3804
rect 19662 3717 19668 3769
rect 19720 3756 19726 3769
rect 19720 3720 92873 3756
rect 19720 3717 19726 3720
rect 19998 3632 20004 3684
rect 20056 3672 20062 3684
rect 20056 3636 92789 3672
rect 20056 3632 20062 3636
rect 20110 3548 20116 3600
rect 20168 3588 20174 3600
rect 20168 3552 92705 3588
rect 20168 3548 20174 3552
rect 21006 3464 21012 3516
rect 21064 3504 21070 3516
rect 21064 3468 92621 3504
rect 21064 3464 21070 3468
rect 21230 3380 21236 3432
rect 21288 3420 21294 3432
rect 21288 3384 92537 3420
rect 21288 3380 21294 3384
rect 21342 3336 21348 3348
rect 21341 3300 21348 3336
rect 21342 3296 21348 3300
rect 21400 3336 21406 3348
rect 21400 3300 92453 3336
rect 21400 3296 21406 3300
rect 21454 3252 21460 3264
rect 21448 3216 21460 3252
rect 21454 3212 21460 3216
rect 21512 3252 21518 3264
rect 21512 3216 92369 3252
rect 21512 3212 21518 3216
rect 29406 3129 29412 3181
rect 29464 3168 29470 3181
rect 29464 3132 92285 3168
rect 29464 3129 29470 3132
rect 29518 3084 29524 3097
rect 29514 3048 29524 3084
rect 29518 3045 29524 3048
rect 29576 3084 29582 3097
rect 29576 3048 92201 3084
rect 29576 3045 29582 3048
rect 29630 3000 29636 3012
rect 29624 2964 29636 3000
rect 29630 2960 29636 2964
rect 29688 3000 29694 3012
rect 29688 2964 92117 3000
rect 29688 2960 29694 2964
rect 29742 2920 29748 2928
rect 29738 2880 29748 2920
rect 29742 2876 29748 2880
rect 29800 2916 29806 2928
rect 29800 2880 92033 2916
rect 29800 2876 29806 2880
rect 21566 2719 21572 2771
rect 21624 2761 21630 2771
rect 83284 2761 83290 2769
rect 21624 2725 83290 2761
rect 21624 2719 21630 2725
rect 83284 2717 83290 2725
rect 83342 2761 83348 2769
rect 83342 2725 83357 2761
rect 83342 2717 83348 2725
rect 21678 2635 21684 2687
rect 21736 2677 21742 2687
rect 83368 2677 83374 2685
rect 21736 2641 83374 2677
rect 21736 2635 21742 2641
rect 83368 2633 83374 2641
rect 83426 2677 83432 2685
rect 83426 2641 83435 2677
rect 83426 2633 83432 2641
rect 21790 2551 21796 2603
rect 21848 2593 21854 2603
rect 83452 2593 83458 2601
rect 21848 2557 83458 2593
rect 21848 2551 21854 2557
rect 83452 2549 83458 2557
rect 83510 2593 83516 2601
rect 83510 2557 83521 2593
rect 83510 2549 83516 2557
rect 21902 2467 21908 2519
rect 21960 2509 21966 2519
rect 83536 2509 83542 2517
rect 21960 2473 83542 2509
rect 21960 2467 21966 2473
rect 83536 2465 83542 2473
rect 83594 2509 83600 2517
rect 83594 2473 83604 2509
rect 83594 2465 83600 2473
rect 83658 2411 83665 2611
rect 31555 2337 31561 2411
rect 31835 2337 83665 2411
rect 83739 2337 83745 2611
rect 91997 2366 92033 2880
rect 92081 2450 92117 2964
rect 92165 2534 92201 3048
rect 92249 2618 92285 3132
rect 92333 2702 92369 3216
rect 92417 2786 92453 3300
rect 92501 2870 92537 3384
rect 92585 2954 92621 3468
rect 92669 3038 92705 3552
rect 92753 3122 92789 3636
rect 92837 3206 92873 3720
rect 92921 3290 92957 3804
rect 93005 3374 93041 3888
rect 93089 3458 93125 3972
rect 93173 3542 93209 4056
rect 93257 3626 93293 4140
rect 93341 3710 93377 4224
rect 93425 3794 93461 4308
rect 93593 3962 93629 4476
rect 93677 4046 93713 4560
rect 93761 4130 93797 4644
rect 93845 4214 93881 4728
rect 93929 4298 93965 4812
rect 94013 4382 94049 4896
rect 94097 4466 94133 4980
rect 94181 4550 94217 5064
rect 94265 4634 94301 5148
rect 94349 4718 94385 5232
rect 94433 4802 94469 5316
rect 94517 4886 94553 5400
rect 94601 4970 94637 5484
rect 94685 5054 94721 5568
rect 290019 5280 290025 5332
rect 290077 5324 290083 5332
rect 543294 5324 543300 5337
rect 290077 5288 543300 5324
rect 290077 5280 290083 5288
rect 543294 5285 543300 5288
rect 543352 5285 543358 5337
rect 289935 5196 289941 5248
rect 289993 5240 289999 5248
rect 544078 5240 544084 5251
rect 289993 5204 544084 5240
rect 289993 5196 289999 5204
rect 544078 5199 544084 5204
rect 544136 5199 544142 5251
rect 289851 5112 289857 5164
rect 289909 5156 289915 5164
rect 544750 5156 544756 5167
rect 289909 5120 544756 5156
rect 289909 5112 289915 5120
rect 544750 5115 544756 5120
rect 544808 5115 544814 5167
rect 286719 5054 286725 5062
rect 94685 5018 286725 5054
rect 286719 5010 286725 5018
rect 286777 5010 286783 5062
rect 289767 5028 289773 5080
rect 289825 5072 289831 5080
rect 545534 5072 545540 5084
rect 289825 5036 545540 5072
rect 289825 5028 289831 5036
rect 545534 5032 545540 5036
rect 545592 5032 545598 5084
rect 286803 4970 286809 4978
rect 94601 4934 286809 4970
rect 286803 4926 286809 4934
rect 286861 4926 286867 4978
rect 289683 4944 289689 4996
rect 289741 4988 289747 4996
rect 549342 4988 549348 5001
rect 289741 4952 549348 4988
rect 289741 4944 289747 4952
rect 549342 4949 549348 4952
rect 549400 4949 549406 5001
rect 286887 4886 286893 4894
rect 94517 4850 286893 4886
rect 286887 4842 286893 4850
rect 286945 4842 286951 4894
rect 289599 4860 289605 4912
rect 289657 4904 289663 4912
rect 549454 4904 549460 4917
rect 289657 4868 549460 4904
rect 289657 4860 289663 4868
rect 549454 4865 549460 4868
rect 549512 4865 549518 4917
rect 286971 4802 286977 4810
rect 94433 4766 286977 4802
rect 286971 4758 286977 4766
rect 287029 4758 287036 4810
rect 289515 4776 289521 4828
rect 289573 4820 289579 4828
rect 549566 4820 549572 4834
rect 289573 4784 549572 4820
rect 289573 4776 289579 4784
rect 549566 4782 549572 4784
rect 549624 4782 549630 4834
rect 247999 4718 248005 4726
rect 94349 4682 248005 4718
rect 247999 4674 248005 4682
rect 248057 4674 248063 4726
rect 289431 4692 289437 4744
rect 289489 4736 289495 4744
rect 549678 4736 549684 4749
rect 289489 4700 549684 4736
rect 289489 4692 289495 4700
rect 549678 4697 549684 4700
rect 549736 4736 549742 4749
rect 549736 4700 549744 4736
rect 549736 4697 549742 4700
rect 248083 4634 248089 4642
rect 94265 4598 248089 4634
rect 248083 4590 248089 4598
rect 248141 4590 248147 4642
rect 289347 4608 289353 4660
rect 289405 4652 289411 4660
rect 549902 4652 549908 4666
rect 289405 4616 549908 4652
rect 289405 4608 289411 4616
rect 549902 4614 549908 4616
rect 549960 4614 549966 4666
rect 248167 4550 248173 4558
rect 94181 4514 248173 4550
rect 248167 4506 248173 4514
rect 248225 4506 248231 4558
rect 289263 4524 289269 4576
rect 289321 4568 289327 4576
rect 550014 4568 550020 4580
rect 289321 4532 550020 4568
rect 289321 4524 289327 4532
rect 550014 4528 550020 4532
rect 550072 4528 550078 4580
rect 248251 4466 248257 4474
rect 94097 4430 248257 4466
rect 248251 4422 248257 4430
rect 248309 4422 248315 4474
rect 289179 4440 289185 4492
rect 289237 4484 289243 4492
rect 550798 4484 550804 4497
rect 289237 4448 550804 4484
rect 289237 4440 289243 4448
rect 550798 4445 550804 4448
rect 550856 4445 550862 4497
rect 287055 4382 287061 4390
rect 94013 4346 287061 4382
rect 287055 4338 287061 4346
rect 287113 4338 287119 4390
rect 289095 4356 289101 4408
rect 289153 4400 289159 4408
rect 550910 4400 550916 4414
rect 289153 4364 550916 4400
rect 289153 4356 289159 4364
rect 550910 4362 550916 4364
rect 550968 4362 550974 4414
rect 287139 4298 287145 4306
rect 93929 4262 287145 4298
rect 287139 4254 287145 4262
rect 287197 4254 287203 4306
rect 289011 4272 289017 4324
rect 289069 4316 289075 4324
rect 551694 4316 551700 4327
rect 289069 4280 551700 4316
rect 289069 4272 289075 4280
rect 551694 4275 551700 4280
rect 551752 4316 551758 4327
rect 551752 4280 551759 4316
rect 551752 4275 551758 4280
rect 287223 4214 287229 4222
rect 93845 4178 287229 4214
rect 287223 4170 287229 4178
rect 287281 4170 287287 4222
rect 288927 4188 288933 4240
rect 288985 4232 288991 4240
rect 551806 4232 551812 4244
rect 288985 4196 551812 4232
rect 288985 4188 288991 4196
rect 551806 4192 551812 4196
rect 551864 4192 551870 4244
rect 287307 4130 287313 4138
rect 93761 4094 287313 4130
rect 287307 4086 287313 4094
rect 287365 4086 287371 4138
rect 288843 4104 288849 4156
rect 288901 4148 288907 4156
rect 551918 4148 551924 4160
rect 288901 4112 551924 4148
rect 288901 4104 288907 4112
rect 551918 4108 551924 4112
rect 551976 4108 551982 4160
rect 248671 4046 248677 4054
rect 93677 4010 248677 4046
rect 248671 4002 248677 4010
rect 248729 4002 248735 4054
rect 288759 4020 288765 4072
rect 288817 4064 288823 4072
rect 552030 4064 552036 4076
rect 288817 4028 552036 4064
rect 288817 4020 288823 4028
rect 552030 4024 552036 4028
rect 552088 4064 552094 4076
rect 552088 4028 552095 4064
rect 552088 4024 552094 4028
rect 248755 3962 248761 3970
rect 93593 3926 248761 3962
rect 248755 3918 248761 3926
rect 248813 3918 248819 3970
rect 288675 3936 288681 3988
rect 288733 3980 288739 3988
rect 552254 3980 552260 3993
rect 288733 3944 552260 3980
rect 288733 3936 288739 3944
rect 552254 3941 552260 3944
rect 552312 3941 552318 3993
rect 288591 3852 288597 3904
rect 288649 3896 288655 3904
rect 552366 3896 552372 3908
rect 288649 3860 552372 3896
rect 288649 3852 288655 3860
rect 552366 3856 552372 3860
rect 552424 3856 552430 3908
rect 248923 3794 248929 3802
rect 93425 3758 248929 3794
rect 248923 3750 248929 3758
rect 248981 3750 248987 3802
rect 288507 3768 288513 3820
rect 288565 3812 288571 3820
rect 553038 3812 553044 3824
rect 288565 3776 553044 3812
rect 288565 3768 288571 3776
rect 553038 3772 553044 3776
rect 553096 3772 553102 3824
rect 249007 3710 249013 3718
rect 93341 3674 249013 3710
rect 249007 3666 249013 3674
rect 249065 3666 249071 3718
rect 288423 3684 288429 3736
rect 288481 3728 288487 3736
rect 553150 3728 553156 3742
rect 288481 3692 553156 3728
rect 288481 3684 288487 3692
rect 553150 3690 553156 3692
rect 553208 3690 553214 3742
rect 287391 3626 287397 3634
rect 93257 3590 287397 3626
rect 287391 3582 287397 3590
rect 287449 3582 287455 3634
rect 288339 3600 288345 3652
rect 288397 3644 288403 3652
rect 553934 3644 553940 3656
rect 288397 3608 553940 3644
rect 288397 3600 288403 3608
rect 553934 3604 553940 3608
rect 553992 3604 553998 3656
rect 287475 3542 287481 3550
rect 93173 3506 287481 3542
rect 287475 3498 287481 3506
rect 287533 3498 287539 3550
rect 288255 3516 288261 3568
rect 288313 3560 288319 3568
rect 554046 3560 554052 3572
rect 288313 3524 554052 3560
rect 288313 3516 288319 3524
rect 554046 3520 554052 3524
rect 554104 3520 554110 3572
rect 287559 3458 287565 3466
rect 93089 3422 287565 3458
rect 287559 3414 287565 3422
rect 287617 3414 287623 3466
rect 288171 3432 288177 3484
rect 288229 3476 288235 3484
rect 554158 3476 554164 3488
rect 288229 3440 554164 3476
rect 288229 3432 288235 3440
rect 554158 3436 554164 3440
rect 554216 3436 554222 3488
rect 287643 3374 287649 3382
rect 93005 3338 287649 3374
rect 287643 3330 287649 3338
rect 287701 3330 287707 3382
rect 288087 3348 288093 3400
rect 288145 3392 288151 3400
rect 554270 3392 554276 3404
rect 288145 3356 554276 3392
rect 288145 3348 288151 3356
rect 554270 3352 554276 3356
rect 554328 3392 554334 3404
rect 554328 3356 554338 3392
rect 554328 3352 554334 3356
rect 249427 3290 249433 3298
rect 92921 3254 249433 3290
rect 249427 3246 249433 3254
rect 249485 3246 249491 3298
rect 288003 3264 288009 3316
rect 288061 3308 288067 3316
rect 554382 3308 554388 3321
rect 288061 3272 554388 3308
rect 288061 3264 288067 3272
rect 554382 3269 554388 3272
rect 554440 3269 554446 3321
rect 249511 3206 249517 3214
rect 92837 3170 249517 3206
rect 249511 3162 249517 3170
rect 249569 3162 249575 3214
rect 287919 3180 287925 3232
rect 287977 3224 287983 3232
rect 554494 3224 554500 3237
rect 287977 3188 554500 3224
rect 287977 3180 287983 3188
rect 554494 3185 554500 3188
rect 554552 3185 554558 3237
rect 249595 3122 249601 3130
rect 92753 3086 249601 3122
rect 249595 3078 249601 3086
rect 249653 3078 249659 3130
rect 287835 3096 287841 3148
rect 287893 3140 287899 3148
rect 554942 3140 554948 3154
rect 287893 3104 554948 3140
rect 287893 3096 287899 3104
rect 554942 3102 554948 3104
rect 555000 3102 555006 3154
rect 249679 3038 249685 3046
rect 92669 3002 249685 3038
rect 249679 2994 249685 3002
rect 249737 2994 249743 3046
rect 287751 3012 287757 3064
rect 287809 3056 287815 3064
rect 555054 3056 555060 3068
rect 287809 3020 555060 3056
rect 287809 3012 287815 3020
rect 555054 3016 555060 3020
rect 555112 3016 555118 3068
rect 249763 2954 249769 2963
rect 92585 2918 249769 2954
rect 249763 2911 249769 2918
rect 249821 2954 249827 2963
rect 249821 2918 249830 2954
rect 249821 2911 249827 2918
rect 363190 2882 363196 2934
rect 363248 2926 363254 2934
rect 490681 2926 490687 2938
rect 363248 2890 490687 2926
rect 363248 2882 363254 2890
rect 249847 2870 249853 2879
rect 92501 2834 249853 2870
rect 249847 2827 249853 2834
rect 249905 2870 249911 2879
rect 490681 2870 490687 2890
rect 490755 2926 490761 2938
rect 534670 2926 534676 2937
rect 490755 2890 534676 2926
rect 490755 2870 490761 2890
rect 534670 2885 534676 2890
rect 534728 2885 534734 2937
rect 249905 2834 249912 2870
rect 467243 2842 467249 2850
rect 249905 2827 249911 2834
rect 467239 2806 467249 2842
rect 467243 2798 467249 2806
rect 467301 2842 467307 2850
rect 534558 2842 534564 2853
rect 467301 2806 534564 2842
rect 467301 2798 467307 2806
rect 534558 2801 534564 2806
rect 534616 2801 534622 2853
rect 249931 2786 249937 2794
rect 92417 2750 249937 2786
rect 249931 2742 249937 2750
rect 249989 2742 249995 2794
rect 467122 2758 467128 2766
rect 467117 2722 467128 2758
rect 467122 2714 467128 2722
rect 467180 2758 467186 2766
rect 534446 2758 534452 2769
rect 467180 2722 534452 2758
rect 467180 2714 467186 2722
rect 534446 2717 534452 2722
rect 534504 2717 534510 2769
rect 250015 2702 250021 2710
rect 92333 2666 250021 2702
rect 250015 2658 250021 2666
rect 250073 2658 250079 2710
rect 467009 2674 467015 2682
rect 467007 2638 467015 2674
rect 467009 2630 467015 2638
rect 467067 2674 467073 2682
rect 534334 2674 534340 2685
rect 467067 2638 534340 2674
rect 467067 2630 467073 2638
rect 534334 2633 534340 2638
rect 534392 2633 534398 2685
rect 286383 2618 286389 2626
rect 92249 2582 286389 2618
rect 286383 2574 286389 2582
rect 286441 2574 286447 2626
rect 466888 2590 466894 2598
rect 466882 2554 466894 2590
rect 466888 2546 466894 2554
rect 466946 2590 466952 2598
rect 534222 2590 534228 2601
rect 466946 2554 534228 2590
rect 466946 2546 466952 2554
rect 534222 2549 534228 2554
rect 534280 2549 534286 2601
rect 286467 2534 286473 2543
rect 92165 2498 286473 2534
rect 286467 2491 286473 2498
rect 286525 2491 286531 2543
rect 469835 2506 469841 2514
rect 469827 2470 469841 2506
rect 469835 2462 469841 2470
rect 469893 2506 469899 2514
rect 534110 2506 534116 2517
rect 469893 2470 534116 2506
rect 469893 2462 469899 2470
rect 534110 2465 534116 2470
rect 534168 2465 534174 2517
rect 286551 2450 286557 2458
rect 92081 2414 286557 2450
rect 286551 2406 286557 2414
rect 286609 2406 286615 2458
rect 469597 2422 469603 2430
rect 469587 2386 469603 2422
rect 469597 2378 469603 2386
rect 469655 2422 469661 2430
rect 533998 2422 534004 2433
rect 469655 2386 534004 2422
rect 469655 2378 469661 2386
rect 533998 2381 534004 2386
rect 534056 2381 534062 2433
rect 286635 2366 286641 2375
rect 91997 2330 286641 2366
rect 286635 2323 286641 2330
rect 286693 2323 286699 2375
rect 469474 2338 469480 2346
rect 469470 2302 469480 2338
rect 469474 2294 469480 2302
rect 469532 2338 469538 2346
rect 533886 2338 533892 2349
rect 469532 2302 533892 2338
rect 469532 2294 469538 2302
rect 533886 2297 533892 2302
rect 533944 2297 533950 2349
rect 22238 2215 22244 2267
rect 22296 2257 22302 2267
rect 22296 2221 232331 2257
rect 472307 2254 472313 2262
rect 22296 2215 22302 2221
rect 472300 2218 472313 2254
rect 472307 2210 472313 2218
rect 472365 2254 472371 2262
rect 533774 2254 533780 2265
rect 472365 2218 533780 2254
rect 472365 2210 472371 2218
rect 533774 2213 533780 2218
rect 533832 2213 533838 2265
rect 22350 2131 22356 2183
rect 22408 2173 22414 2183
rect 194587 2173 194593 2181
rect 22408 2137 194593 2173
rect 22408 2131 22414 2137
rect 194587 2129 194593 2137
rect 194645 2173 194651 2181
rect 194645 2137 194682 2173
rect 472431 2170 472437 2178
rect 194645 2129 194651 2137
rect 472422 2134 472437 2170
rect 472431 2126 472437 2134
rect 472489 2170 472495 2178
rect 533662 2170 533668 2181
rect 472489 2134 533668 2170
rect 472489 2126 472495 2134
rect 533662 2129 533668 2134
rect 533720 2129 533726 2181
rect 22462 2047 22468 2099
rect 22520 2089 22526 2099
rect 197070 2089 197076 2096
rect 22520 2053 197076 2089
rect 22520 2047 22526 2053
rect 197070 2044 197076 2053
rect 197128 2044 197134 2096
rect 472185 2086 472191 2094
rect 472180 2050 472191 2086
rect 472185 2042 472191 2050
rect 472243 2086 472249 2094
rect 533550 2086 533556 2097
rect 472243 2050 533556 2086
rect 472243 2042 472249 2050
rect 533550 2045 533556 2050
rect 533608 2045 533614 2097
rect 22574 1963 22580 2015
rect 22632 2005 22638 2015
rect 22632 1996 174822 2005
rect 472067 2002 472073 2010
rect 22632 1969 174729 1996
rect 174781 1969 174822 1996
rect 22632 1963 22638 1969
rect 472056 1966 472073 2002
rect 472067 1958 472073 1966
rect 472125 2002 472131 2010
rect 533438 2002 533444 2013
rect 472125 1966 533444 2002
rect 472125 1958 472131 1966
rect 533438 1961 533444 1966
rect 533496 1961 533502 2013
rect 22686 1879 22692 1931
rect 22744 1921 22750 1931
rect 135648 1921 135654 1929
rect 22744 1885 135654 1921
rect 22744 1879 22750 1885
rect 135648 1877 135654 1885
rect 135706 1921 135712 1929
rect 135706 1885 135739 1921
rect 474901 1918 474907 1926
rect 135706 1877 135712 1885
rect 474895 1882 474907 1918
rect 474901 1874 474907 1882
rect 474959 1918 474965 1926
rect 533326 1918 533332 1929
rect 474959 1882 533332 1918
rect 474959 1874 474965 1882
rect 533326 1877 533332 1882
rect 533384 1877 533390 1929
rect 22798 1795 22804 1847
rect 22856 1837 22862 1847
rect 138104 1837 138110 1844
rect 22856 1801 138110 1837
rect 22856 1795 22862 1801
rect 138104 1792 138110 1801
rect 138162 1837 138168 1844
rect 138162 1801 138174 1837
rect 475022 1834 475028 1842
rect 138162 1792 138168 1801
rect 475020 1798 475028 1834
rect 475022 1790 475028 1798
rect 475080 1834 475086 1842
rect 533214 1834 533220 1845
rect 475080 1798 533220 1834
rect 475080 1790 475086 1798
rect 533214 1793 533220 1798
rect 533272 1793 533278 1845
rect 22910 1711 22916 1763
rect 22968 1753 22974 1763
rect 189211 1753 189217 1761
rect 22968 1717 189217 1753
rect 22968 1711 22974 1717
rect 189211 1709 189217 1717
rect 189269 1709 189275 1761
rect 474779 1750 474785 1758
rect 474769 1714 474785 1750
rect 474779 1706 474785 1714
rect 474837 1750 474843 1758
rect 533102 1750 533108 1761
rect 474837 1714 533108 1750
rect 474837 1706 474843 1714
rect 533102 1709 533108 1714
rect 533160 1709 533166 1761
rect 20443 1625 20449 1677
rect 20501 1669 20507 1677
rect 273394 1669 273400 1678
rect 20501 1633 273400 1669
rect 20501 1625 20507 1633
rect 273394 1626 273400 1633
rect 273452 1669 273458 1678
rect 273452 1633 273459 1669
rect 474658 1666 474664 1674
rect 273452 1626 273458 1633
rect 474653 1630 474664 1666
rect 474658 1622 474664 1630
rect 474716 1666 474722 1674
rect 532990 1666 532996 1677
rect 474716 1630 532996 1666
rect 474716 1622 474722 1630
rect 532990 1625 532996 1630
rect 533048 1625 533054 1677
rect 20555 1541 20561 1593
rect 20613 1585 20619 1593
rect 273478 1585 273484 1594
rect 20613 1549 273484 1585
rect 20613 1541 20619 1549
rect 273478 1542 273484 1549
rect 273536 1585 273542 1594
rect 273536 1549 273545 1585
rect 477492 1582 477498 1590
rect 273536 1542 273542 1549
rect 477482 1546 477498 1582
rect 477492 1538 477498 1546
rect 477550 1582 477556 1590
rect 532878 1582 532884 1593
rect 477550 1546 532884 1582
rect 477550 1538 477556 1546
rect 532878 1541 532884 1546
rect 532936 1541 532942 1593
rect 20672 1457 20678 1509
rect 20730 1501 20736 1509
rect 273562 1501 273568 1510
rect 20730 1465 273568 1501
rect 20730 1457 20736 1465
rect 273562 1458 273568 1465
rect 273620 1501 273626 1510
rect 273620 1465 273632 1501
rect 469716 1498 469722 1506
rect 273620 1458 273626 1465
rect 469712 1462 469722 1498
rect 469716 1454 469722 1462
rect 469774 1498 469780 1506
rect 532766 1498 532772 1509
rect 469774 1462 532772 1498
rect 469774 1454 469780 1462
rect 532766 1457 532772 1462
rect 532824 1457 532830 1509
rect 20784 1373 20790 1425
rect 20842 1417 20848 1425
rect 273646 1417 273652 1426
rect 20842 1381 273652 1417
rect 20842 1373 20848 1381
rect 273646 1374 273652 1381
rect 273704 1417 273710 1426
rect 482804 1422 482856 1428
rect 273704 1381 273713 1417
rect 273704 1374 273710 1381
rect 482790 1378 482804 1414
rect 532654 1414 532660 1425
rect 482856 1378 532660 1414
rect 532654 1373 532660 1378
rect 532712 1373 532718 1425
rect 482804 1364 482856 1370
rect 482555 1330 482561 1338
rect 482549 1294 482561 1330
rect 482555 1286 482561 1294
rect 482613 1330 482619 1338
rect 532542 1330 532548 1341
rect 482613 1294 532548 1330
rect 482613 1286 482619 1294
rect 532542 1289 532548 1294
rect 532600 1289 532606 1341
rect 477608 1246 477614 1254
rect 477602 1210 477614 1246
rect 477608 1202 477614 1210
rect 477666 1246 477672 1254
rect 532430 1246 532436 1257
rect 477666 1210 532436 1246
rect 477666 1202 477672 1210
rect 532430 1205 532436 1210
rect 532488 1205 532494 1257
rect 477373 1162 477379 1170
rect 477367 1126 477379 1162
rect 477373 1118 477379 1126
rect 477431 1162 477437 1170
rect 532318 1162 532324 1173
rect 477431 1126 532324 1162
rect 477431 1118 477437 1126
rect 532318 1121 532324 1126
rect 532376 1121 532382 1173
rect 477252 1034 477258 1086
rect 477310 1078 477316 1086
rect 532206 1078 532212 1089
rect 477310 1042 532212 1078
rect 477310 1034 477316 1042
rect 532206 1037 532212 1042
rect 532264 1037 532270 1089
rect 482439 994 482445 1002
rect 482433 958 482445 994
rect 482439 950 482445 958
rect 482497 994 482503 1002
rect 532094 994 532100 1005
rect 482497 958 532100 994
rect 482497 950 482503 958
rect 532094 953 532100 958
rect 532152 953 532158 1005
rect 482679 910 482685 918
rect 482676 874 482685 910
rect 482679 866 482685 874
rect 482737 910 482743 918
rect 531982 910 531988 921
rect 482737 874 531988 910
rect 482737 866 482743 874
rect 531982 869 531988 874
rect 532040 869 532046 921
rect 480085 826 480091 834
rect 480081 790 480091 826
rect 480085 782 480091 790
rect 480143 826 480149 834
rect 531870 826 531876 837
rect 480143 790 531876 826
rect 480143 782 480149 790
rect 531870 785 531876 790
rect 531928 785 531934 837
rect 480201 742 480207 750
rect 480194 706 480207 742
rect 480201 698 480207 706
rect 480259 742 480265 750
rect 531758 742 531764 753
rect 480259 706 531764 742
rect 480259 698 480265 706
rect 531758 701 531764 706
rect 531816 701 531822 753
rect 479960 658 479966 666
rect 479949 622 479966 658
rect 479960 614 479966 622
rect 480018 658 480024 666
rect 531646 658 531652 669
rect 480018 622 531652 658
rect 480018 614 480024 622
rect 531646 617 531652 622
rect 531704 617 531710 669
rect 479841 574 479847 582
rect 479834 538 479847 574
rect 479841 530 479847 538
rect 479899 574 479905 582
rect 531534 574 531540 585
rect 479899 538 531540 574
rect 479899 530 479905 538
rect 531534 533 531540 538
rect 531592 533 531598 585
rect 363271 490 363277 498
rect 363264 454 363277 490
rect 363271 446 363277 454
rect 363329 490 363335 498
rect 531422 490 531428 501
rect 363329 454 531428 490
rect 363329 446 363335 454
rect 531422 449 531428 454
rect 531480 449 531486 501
<< via1 >>
rect 504656 110336 504708 110388
rect 504536 110216 504588 110268
rect 504896 110096 504948 110148
rect 504774 109976 504826 110028
rect 498988 109856 499040 109908
rect 498876 109736 498928 109788
rect 498746 109616 498798 109668
rect 498626 109496 498678 109548
rect 321596 109376 321648 109428
rect 321718 109256 321770 109308
rect 321350 109136 321402 109188
rect 91305 109017 91357 109069
rect 321468 109016 321520 109068
rect 91182 108945 91234 108997
rect 91052 108873 91104 108925
rect 315446 108896 315498 108948
rect 90936 108801 90988 108853
rect 96965 108729 97017 108781
rect 315558 108776 315610 108828
rect 96846 108657 96898 108709
rect 315678 108656 315730 108708
rect 97208 108585 97260 108637
rect 97084 108513 97136 108565
rect 315804 108536 315856 108588
rect 267209 108437 267261 108489
rect 267089 108365 267141 108417
rect 266964 108293 267016 108345
rect 266840 108221 266892 108273
rect 272872 108149 272924 108201
rect 272747 108077 272799 108129
rect 266840 107819 266892 107871
rect 266963 107816 267015 107868
rect 90936 107677 90988 107729
rect 91059 107686 91111 107738
rect 267085 107802 267137 107854
rect 267210 107812 267262 107864
rect 272747 107840 272799 107892
rect 272872 107849 272924 107901
rect 91182 107670 91234 107722
rect 91298 107677 91350 107729
rect 96846 107659 96898 107711
rect 96965 107647 97017 107699
rect 97084 107668 97136 107720
rect 321350 107886 321402 107938
rect 321468 107886 321520 107938
rect 321596 107896 321648 107948
rect 321718 107898 321770 107950
rect 315446 107710 315498 107762
rect 315556 107720 315608 107772
rect 315678 107734 315730 107786
rect 315804 107734 315856 107786
rect 97208 107647 97260 107699
rect 498626 107818 498678 107870
rect 498746 107806 498798 107858
rect 498876 107808 498928 107860
rect 498988 107806 499040 107858
rect 504536 107808 504588 107860
rect 504656 107818 504708 107870
rect 504774 107830 504826 107882
rect 504896 107828 504948 107880
rect 509025 107274 509105 107354
rect 508926 104866 509006 104946
rect 48440 104470 48520 104550
rect 45400 102542 45452 102594
rect 45316 102458 45368 102510
rect 45232 102374 45284 102426
rect 45148 102291 45200 102343
rect 45064 102206 45116 102258
rect 44980 102121 45032 102173
rect 46912 102039 46964 102091
rect 48330 102070 48410 102150
rect 46828 101955 46880 102007
rect 46744 101870 46796 101922
rect 46660 101786 46712 101838
rect 46576 101703 46628 101755
rect 46492 101620 46544 101672
rect 48230 99700 48310 99780
rect 48120 97300 48200 97380
rect 47416 96676 47468 96728
rect 47332 96592 47384 96644
rect 47248 96509 47300 96561
rect 47164 96425 47216 96477
rect 47080 96339 47132 96391
rect 46996 96258 47048 96310
rect 46408 96174 46460 96226
rect 46324 96089 46376 96141
rect 46240 96006 46292 96058
rect 46156 95920 46208 95972
rect 46072 95840 46124 95892
rect 45988 95752 46040 95804
rect 48014 94900 48094 94980
rect 45904 90809 45956 90861
rect 45820 90728 45872 90780
rect 45736 90643 45788 90695
rect 45652 90559 45704 90611
rect 45568 90475 45620 90527
rect 45484 90391 45536 90443
rect 47500 90308 47552 90360
rect 47920 90222 47972 90274
rect 47836 90138 47888 90190
rect 47752 90054 47804 90106
rect 47668 89970 47720 90022
rect 47584 89886 47636 89938
rect 10148 84052 10200 84104
rect 10260 83926 10312 83978
rect 10372 83804 10424 83856
rect 10484 83689 10536 83741
rect 9924 78142 9976 78194
rect 10036 78013 10088 78065
rect 9700 77901 9752 77953
rect 9812 77777 9864 77829
rect 28889 77323 28941 77375
rect 28973 77239 29025 77291
rect 29057 77155 29109 77207
rect 286469 102999 286531 103061
rect 286389 102716 286441 102768
rect 508830 102468 508910 102548
rect 287314 101124 287366 101176
rect 287230 101040 287282 101092
rect 287733 100957 287785 101009
rect 287817 100875 287869 100927
rect 287061 100789 287113 100841
rect 287145 100704 287197 100756
rect 508740 100088 508820 100168
rect 508642 97672 508722 97752
rect 286893 93253 286945 93305
rect 286977 93172 287029 93224
rect 287480 93086 287532 93138
rect 287398 93002 287450 93054
rect 287565 92917 287617 92969
rect 287649 92836 287701 92888
rect 48550 92517 48602 92569
rect 48532 90100 48612 90180
rect 29141 77071 29193 77123
rect 48365 87694 48417 87746
rect 48261 85318 48313 85370
rect 29225 76987 29277 77039
rect 48157 82910 48213 82966
rect 29309 76903 29361 76955
rect 29393 76819 29445 76871
rect 29477 76735 29529 76787
rect 29561 76651 29613 76703
rect 388908 90725 390258 90856
rect 434187 90780 435612 90895
rect 198858 90469 200372 90609
rect 154585 90232 156040 90355
rect 196222 89834 196274 89886
rect 158300 89591 158352 89643
rect 388995 89177 390345 89308
rect 198845 88930 200359 89070
rect 154673 88696 156003 88824
rect 29645 76567 29697 76619
rect 286636 86946 286696 87006
rect 286557 86650 286609 86702
rect 286810 85048 286862 85100
rect 286725 84964 286777 85016
rect 287146 84880 287198 84932
rect 287062 84796 287114 84848
rect 289605 84712 289657 84764
rect 289689 84627 289741 84679
rect 287985 83284 288037 83336
rect 289017 83286 289069 83338
rect 287901 83200 287953 83252
rect 288933 83202 288985 83254
rect 287817 83116 287869 83168
rect 288849 83118 288901 83170
rect 287733 83032 287785 83084
rect 288765 83034 288817 83086
rect 287313 82949 287365 83001
rect 288345 82948 288397 83000
rect 287229 82865 287281 82917
rect 288261 82864 288313 82916
rect 286977 82782 287029 82834
rect 288177 82780 288229 82832
rect 286893 82698 286945 82750
rect 288093 82696 288145 82748
rect 48765 80907 49066 81227
rect 48765 79677 49066 79997
rect 29729 76483 29781 76535
rect 163169 77986 163221 78038
rect 29813 76399 29865 76451
rect 158300 77903 158352 77955
rect 94230 77783 94282 77835
rect 94314 77699 94366 77751
rect 94398 77615 94450 77667
rect 94482 77531 94534 77583
rect 94566 77447 94618 77499
rect 94650 77363 94702 77415
rect 94734 77279 94786 77331
rect 94818 77195 94870 77247
rect 94902 77111 94954 77163
rect 94986 77027 95038 77079
rect 95070 76943 95122 76995
rect 95154 76859 95206 76911
rect 95238 76775 95290 76827
rect 95322 76691 95374 76743
rect 95406 76607 95458 76659
rect 95490 76523 95542 76575
rect 434639 89231 435961 89367
rect 507538 79888 507590 79940
rect 507622 79805 507674 79857
rect 507707 79721 507759 79773
rect 507791 79636 507843 79688
rect 507875 79552 507927 79604
rect 507959 79469 508011 79521
rect 508043 79383 508095 79435
rect 508127 79300 508179 79352
rect 507454 79217 507506 79269
rect 507370 79133 507422 79185
rect 507286 79049 507338 79101
rect 507202 78965 507254 79017
rect 507118 78881 507170 78933
rect 507034 78797 507086 78849
rect 506950 78713 507002 78765
rect 506866 78629 506918 78681
rect 509485 95282 509565 95362
rect 509398 92892 509478 92972
rect 509303 90482 509383 90562
rect 509230 88119 509282 88171
rect 509147 85702 509199 85754
rect 568824 88934 568876 88986
rect 568936 88820 568988 88872
rect 569048 88700 569100 88752
rect 569160 88566 569212 88618
rect 509759 83681 510920 83844
rect 569272 83022 569324 83074
rect 569384 82904 569436 82956
rect 569496 82784 569548 82836
rect 509771 82541 510932 82704
rect 569608 82670 569660 82722
rect 376248 78324 376300 78376
rect 510402 78402 510454 78454
rect 380666 78227 380718 78279
rect 510318 78318 510370 78370
rect 458770 78230 458822 78282
rect 510234 78234 510286 78286
rect 385200 78145 385252 78197
rect 510150 78150 510202 78202
rect 482242 78066 482294 78118
rect 510066 78066 510118 78118
rect 191486 77986 191538 78038
rect 196222 77986 196274 78038
rect 445190 77988 445242 78040
rect 509982 77982 510034 78034
rect 440456 77896 440508 77948
rect 509898 77898 509950 77950
rect 454384 77812 454436 77864
rect 509814 77814 509866 77866
rect 435838 77724 435890 77776
rect 509730 77730 509782 77782
rect 477526 77644 477578 77696
rect 509646 77646 509698 77698
rect 463586 77564 463638 77616
rect 509562 77562 509614 77614
rect 486858 77480 486910 77532
rect 509478 77478 509530 77530
rect 468232 77392 468284 77444
rect 509394 77394 509446 77446
rect 491474 77312 491526 77364
rect 509310 77310 509362 77362
rect 528470 78258 528522 78310
rect 528386 78174 528438 78226
rect 528302 78090 528354 78142
rect 528218 78006 528270 78058
rect 528134 77922 528186 77974
rect 528050 77838 528102 77890
rect 527966 77754 528018 77806
rect 527882 77670 527934 77722
rect 527798 77586 527850 77638
rect 527714 77502 527766 77554
rect 528638 77323 528690 77375
rect 289437 77178 289489 77230
rect 528557 77227 528609 77279
rect 289521 77094 289573 77146
rect 286978 77010 287030 77062
rect 286894 76926 286946 76978
rect 287312 76842 287364 76894
rect 287229 76758 287281 76810
rect 34596 76025 34648 76077
rect 231378 76024 231430 76076
rect 34680 75941 34732 75993
rect 199064 75946 199116 75998
rect 34764 75857 34816 75909
rect 219892 75860 219944 75912
rect 34848 75773 34900 75825
rect 203482 75779 203534 75831
rect 34932 75689 34984 75741
rect 208016 75691 208068 75743
rect 35016 75605 35068 75657
rect 235894 75608 235946 75660
rect 35100 75521 35152 75573
rect 152454 75528 152506 75580
rect 35184 75437 35236 75489
rect 224408 75438 224460 75490
rect 35268 75353 35320 75405
rect 147920 75356 147972 75408
rect 35352 75269 35404 75321
rect 143502 75269 143554 75321
rect 35436 75185 35488 75237
rect 240410 75183 240462 75235
rect 35520 75101 35572 75153
rect 215376 75100 215428 75152
rect 527414 77140 527466 77192
rect 526838 77056 526890 77108
rect 526478 76972 526530 77024
rect 525326 76890 525378 76942
rect 527198 76804 527250 76856
rect 527054 76720 527106 76772
rect 526694 76636 526746 76688
rect 525758 76552 525810 76604
rect 527342 76468 527394 76520
rect 526766 76384 526818 76436
rect 526406 76300 526458 76352
rect 525254 76216 525306 76268
rect 527126 76134 527178 76186
rect 526982 76048 527034 76100
rect 526622 75964 526674 76016
rect 525686 75882 525738 75934
rect 524822 75796 524874 75848
rect 525038 75712 525090 75764
rect 526334 75628 526386 75680
rect 525614 75544 525666 75596
rect 526910 75462 526962 75514
rect 525398 75376 525450 75428
rect 526550 75290 526602 75342
rect 524174 65774 524226 65826
rect 523670 65690 523722 65742
rect 525830 65606 525882 65658
rect 524462 65522 524514 65574
rect 523958 65438 524010 65490
rect 526118 65358 526170 65410
rect 527270 65270 527322 65322
rect 524246 65186 524298 65238
rect 523742 65104 523794 65156
rect 525902 65020 525954 65072
rect 525470 64934 525522 64986
rect 524678 64850 524730 64902
rect 524534 64768 524586 64820
rect 524030 64682 524082 64734
rect 526190 64598 526242 64650
rect 525110 64514 525162 64566
rect 524894 64432 524946 64484
rect 524318 64346 524370 64398
rect 523814 64262 523866 64314
rect 525974 64178 526026 64230
rect 525542 64094 525594 64146
rect 524750 64010 524802 64062
rect 524606 63926 524658 63978
rect 524102 63842 524154 63894
rect 526262 63758 526314 63810
rect 525182 63674 525234 63726
rect 524966 63590 525018 63642
rect 524390 63506 524442 63558
rect 523886 63422 523938 63474
rect 526046 63338 526098 63390
rect 385990 63241 386042 63293
rect 544430 63240 544482 63292
rect 416042 63158 416094 63210
rect 480551 63156 480603 63208
rect 544346 63156 544398 63208
rect 415958 63074 416010 63126
rect 480635 63072 480687 63124
rect 544262 63072 544314 63124
rect 415874 62990 415926 63042
rect 480719 62988 480771 63040
rect 544178 62988 544230 63040
rect 415790 62905 415842 62957
rect 480803 62904 480855 62956
rect 544094 62904 544146 62956
rect 480887 62820 480939 62872
rect 544010 62820 544062 62872
rect 480971 62736 481023 62788
rect 543926 62736 543978 62788
rect 481055 62652 481107 62704
rect 543842 62652 543894 62704
rect 481139 62568 481191 62620
rect 543758 62568 543810 62620
rect 481223 62484 481275 62536
rect 543674 62484 543726 62536
rect 481307 62400 481359 62452
rect 543590 62400 543642 62452
rect 481391 62316 481443 62368
rect 543506 62316 543558 62368
rect 481475 62232 481527 62284
rect 543422 62232 543474 62284
rect 374013 62170 374065 62222
rect 374135 62086 374187 62138
rect 83665 61744 83739 61969
rect 84254 61906 84306 61958
rect 292066 61889 292118 61941
rect 292150 61805 292202 61857
rect 340623 61722 340675 61774
rect 340539 61638 340591 61690
rect 289941 61451 289993 61503
rect 290025 61370 290077 61422
rect 183998 59273 185192 59797
rect 83288 58763 83340 58815
rect 30174 57165 30226 57217
rect 76404 57165 76456 57217
rect 30005 57081 30057 57133
rect 70609 57081 70661 57133
rect 30089 56997 30141 57049
rect 69968 56997 70020 57049
rect 31013 56913 31065 56965
rect 67378 56913 67430 56965
rect 30846 56829 30898 56881
rect 64933 56829 64985 56881
rect 9252 55843 9304 55895
rect 9364 55716 9416 55768
rect 9476 55611 9528 55663
rect 9589 55493 9641 55545
rect 289773 61289 289825 61341
rect 289860 61205 289912 61257
rect 340455 61554 340507 61606
rect 292320 61471 292372 61523
rect 292404 61385 292456 61437
rect 292485 61301 292537 61353
rect 292236 61218 292288 61270
rect 374254 61133 374306 61185
rect 341058 61025 341158 61125
rect 391306 60956 391358 61008
rect 481559 62148 481611 62200
rect 543338 62148 543390 62200
rect 481643 62064 481695 62116
rect 543254 62064 543306 62116
rect 481727 61980 481779 62032
rect 543170 61980 543222 62032
rect 481811 61896 481863 61948
rect 543086 61896 543138 61948
rect 415706 61812 415758 61864
rect 543002 61812 543054 61864
rect 542918 61728 542970 61780
rect 542834 61644 542886 61696
rect 429774 61522 430184 61588
rect 430758 61564 431270 61622
rect 430717 61470 430769 61522
rect 522215 61471 522267 61523
rect 430800 61386 430852 61438
rect 522131 61386 522183 61438
rect 522319 61395 522371 61607
rect 542750 61302 542802 61354
rect 542666 61218 542718 61270
rect 542582 61134 542634 61186
rect 542498 61050 542550 61102
rect 485628 60966 485680 61018
rect 519080 60966 519132 61018
rect 542414 60966 542466 61018
rect 485712 60882 485764 60934
rect 518996 60882 519048 60934
rect 542330 60882 542382 60934
rect 485794 60798 485846 60850
rect 518912 60798 518964 60850
rect 542246 60798 542298 60850
rect 485882 60714 485934 60766
rect 518828 60714 518880 60766
rect 542162 60714 542214 60766
rect 485968 60630 486020 60682
rect 518744 60630 518796 60682
rect 542078 60630 542130 60682
rect 481937 60547 481989 60599
rect 486046 60546 486098 60598
rect 518660 60546 518712 60598
rect 541994 60546 542046 60598
rect 486136 60462 486188 60514
rect 518576 60462 518628 60514
rect 541910 60462 541962 60514
rect 561010 60460 561062 60512
rect 486216 60378 486268 60430
rect 518492 60378 518544 60430
rect 541826 60378 541878 60430
rect 422513 60294 422565 60346
rect 486298 60294 486350 60346
rect 518408 60294 518460 60346
rect 541742 60294 541794 60346
rect 486382 60210 486434 60262
rect 518324 60210 518376 60262
rect 541658 60210 541710 60262
rect 486468 60126 486520 60178
rect 518240 60126 518292 60178
rect 541574 60126 541626 60178
rect 406725 59616 407761 59916
rect 342790 58606 342918 59266
rect 343302 58606 343430 59266
rect 343814 58606 343942 59266
rect 344326 58606 344454 59266
rect 344838 58606 344966 59266
rect 345350 58606 345478 59266
rect 345862 58606 345990 59266
rect 346374 58606 346502 59266
rect 346886 58606 347014 59266
rect 347398 58606 347526 59266
rect 348422 58606 348550 59266
rect 348934 58606 349062 59266
rect 349446 58606 349574 59266
rect 349958 58606 350086 59266
rect 350470 58606 350598 59266
rect 350982 58606 351110 59266
rect 351494 58606 351622 59266
rect 352180 58638 353960 59225
rect 288010 56759 288062 56811
rect 288510 56675 288562 56727
rect 289188 56591 289240 56643
rect 354362 54424 354414 54476
rect 186242 53968 186294 54020
rect 83370 52496 83422 52548
rect 186566 52384 187774 52604
rect 249601 52115 249653 52167
rect 287836 52126 287888 52178
rect 288684 52042 288736 52094
rect 248173 51956 248225 52008
rect 289356 51958 289408 52010
rect 248677 51866 248729 51918
rect 249433 51786 249485 51838
rect 248929 51661 248981 51713
rect 250547 51665 250599 51717
rect 241594 51575 241646 51627
rect 249769 51575 249821 51627
rect 241895 51432 241947 51484
rect 249853 51436 249905 51488
rect 241510 51305 241562 51357
rect 249937 51302 249989 51354
rect 246019 51140 246071 51192
rect 248007 51140 248059 51192
rect 241176 51022 241228 51074
rect 250022 51022 250074 51074
rect 9028 49934 9080 49986
rect 9140 49824 9192 49876
rect 522299 49862 522351 50114
rect 354284 49792 354336 49844
rect 522215 49778 522267 49830
rect 540164 49784 540216 49836
rect 8804 49697 8856 49749
rect 522131 49693 522183 49745
rect 540052 49699 540104 49751
rect 540273 49693 540332 49920
rect 8916 49581 8968 49633
rect 374013 48873 374065 48925
rect 374135 48768 374187 48820
rect 374254 48664 374306 48716
rect 248082 47493 248134 47545
rect 287929 47493 287981 47545
rect 422514 47518 422566 47570
rect 249009 47409 249061 47461
rect 288428 47409 288480 47461
rect 249687 47325 249739 47377
rect 289103 47325 289155 47377
rect 562759 60236 564261 60665
rect 561926 60176 561978 60228
rect 561250 60082 561302 60134
rect 562408 60094 562460 60146
rect 562048 60010 562100 60062
rect 562646 59938 562698 59990
rect 564801 59866 564853 59918
rect 561128 59794 561180 59846
rect 561690 59722 561742 59774
rect 562168 59650 562220 59702
rect 562528 59578 562580 59630
rect 565210 58543 566611 58968
rect 568608 54618 568660 54670
rect 568724 54498 568776 54550
rect 567712 54368 567764 54420
rect 567824 54260 567876 54312
rect 567488 48710 567540 48762
rect 567600 48596 567652 48648
rect 567264 48470 567316 48522
rect 567376 48346 567428 48398
rect 561570 48056 561622 48108
rect 562288 47976 562340 48028
rect 562770 47896 562822 47948
rect 562886 47816 562938 47868
rect 560962 47656 561014 47708
rect 561088 47542 561140 47594
rect 560722 47416 560774 47468
rect 560844 47296 560896 47348
rect 420803 47023 421743 47148
rect 567936 47124 567988 47176
rect 83460 46845 83512 46897
rect 403905 46006 404057 46464
rect 404206 46000 404358 46458
rect 420789 46034 421670 46173
rect 415706 45844 415758 45896
rect 415790 45753 415842 45805
rect 415874 45667 415926 45719
rect 353772 45160 353824 45212
rect 391672 45018 392309 45630
rect 402906 45570 402958 45622
rect 415958 45569 416010 45621
rect 402908 45463 402960 45515
rect 416042 45462 416094 45514
rect 452727 44712 452779 44764
rect 480551 44709 480603 44761
rect 446720 44628 446772 44680
rect 480635 44625 480687 44677
rect 452565 44544 452617 44596
rect 480719 44541 480771 44593
rect 446884 44460 446936 44512
rect 480803 44457 480855 44509
rect 452405 44376 452457 44428
rect 480887 44373 480939 44425
rect 447043 44292 447095 44344
rect 480971 44289 481023 44341
rect 452243 44208 452295 44260
rect 481055 44205 481107 44257
rect 447207 44124 447259 44176
rect 481139 44121 481191 44173
rect 452088 44040 452140 44092
rect 481223 44037 481275 44089
rect 447365 43956 447417 44008
rect 481307 43953 481359 44005
rect 451920 43872 451972 43924
rect 481391 43869 481443 43921
rect 447524 43788 447576 43840
rect 481475 43785 481527 43837
rect 451765 43704 451817 43756
rect 481559 43701 481611 43753
rect 447688 43620 447740 43672
rect 481643 43617 481695 43669
rect 451603 43536 451655 43588
rect 481727 43533 481779 43585
rect 447846 43452 447898 43504
rect 481811 43449 481863 43501
rect 248259 42860 248311 42912
rect 287764 42860 287816 42912
rect 248758 42776 248810 42828
rect 288594 42776 288646 42828
rect 249515 42692 249567 42744
rect 289271 42692 289323 42744
rect 353188 42608 353240 42660
rect 353272 42324 353324 42376
rect 8356 41856 8408 41908
rect 452125 41808 459416 42875
rect 8468 41731 8520 41783
rect 8580 41606 8632 41658
rect 473111 41785 480402 42852
rect 8692 41491 8744 41543
rect 568048 47000 568100 47052
rect 567040 41384 567092 41436
rect 567152 41262 567204 41314
rect 566816 41130 566868 41182
rect 566928 41026 566980 41078
rect 83546 40578 83598 40630
rect 353696 39374 353748 39426
rect 353020 37630 353072 37682
rect 353104 37342 353156 37394
rect 7908 35945 7960 35997
rect 8020 35824 8072 35876
rect 8132 35706 8184 35758
rect 8244 35581 8296 35633
rect 566592 35478 566644 35530
rect 566704 35350 566756 35402
rect 566368 35244 566420 35296
rect 566480 35104 566532 35156
rect 568384 34704 568436 34756
rect 568496 34560 568548 34612
rect 353858 34378 353910 34430
rect 568160 33468 568212 33520
rect 352852 32666 352904 32718
rect 352936 32376 352988 32428
rect 273484 31262 273536 31314
rect 273400 31141 273452 31193
rect 353944 29432 353996 29484
rect 233042 28332 233094 28384
rect 173952 27872 174004 27924
rect 568272 33374 568324 33426
rect 566144 27986 566196 28038
rect 566256 27878 566308 27930
rect 565920 27764 565972 27816
rect 7460 27666 7512 27718
rect 352684 27684 352736 27736
rect 566032 27634 566084 27686
rect 7572 27540 7624 27592
rect 7684 27413 7736 27465
rect 352768 27380 352820 27432
rect 7796 27290 7848 27342
rect 257258 24982 257372 26004
rect 273652 25355 273704 25407
rect 273568 25234 273620 25286
rect 354026 24470 354078 24522
rect 353524 22698 353576 22750
rect 353608 22404 353660 22456
rect 7236 21744 7288 21796
rect 431923 21785 438850 22602
rect 7348 21625 7400 21677
rect 473177 21637 478353 22662
rect 569280 22092 569332 22144
rect 7012 21512 7064 21564
rect 569392 21970 569444 22022
rect 568832 21838 568884 21890
rect 568944 21736 568996 21788
rect 569056 21618 569108 21670
rect 569168 21510 569220 21562
rect 7124 21391 7176 21443
rect 467480 21247 467532 21299
rect 530452 21297 530504 21349
rect 540943 21297 540995 21349
rect 465398 21161 465450 21213
rect 465066 21076 465118 21128
rect 464770 20995 464822 21047
rect 464469 20909 464521 20961
rect 354110 19566 354162 19618
rect 354194 19446 354246 19498
rect 354364 19304 354416 19356
rect 482496 19944 482548 19996
rect 354280 19220 354332 19272
rect 482412 19860 482464 19912
rect 354196 19136 354248 19188
rect 482328 19776 482380 19828
rect 294545 16433 295010 19081
rect 354112 19052 354164 19104
rect 482244 19692 482296 19744
rect 354028 18968 354080 19020
rect 482160 19608 482212 19660
rect 353944 18884 353996 18936
rect 482076 19524 482128 19576
rect 353860 18800 353912 18852
rect 481992 19440 482044 19492
rect 353776 18716 353828 18768
rect 481908 19356 481960 19408
rect 353692 18632 353744 18684
rect 481824 19272 481876 19324
rect 353608 18548 353660 18600
rect 481740 19188 481792 19240
rect 353524 18464 353576 18516
rect 481656 19104 481708 19156
rect 353392 18380 353444 18432
rect 481572 19020 481624 19072
rect 352572 18296 352624 18348
rect 481488 18936 481540 18988
rect 353272 18212 353324 18264
rect 481404 18852 481456 18904
rect 353188 18128 353240 18180
rect 481320 18768 481372 18820
rect 353104 18044 353156 18096
rect 481236 18684 481288 18736
rect 353020 17960 353072 18012
rect 481152 18600 481204 18652
rect 352936 17876 352988 17928
rect 481068 18516 481120 18568
rect 352852 17792 352904 17844
rect 480984 18432 481036 18484
rect 352572 17732 352624 17784
rect 352768 17708 352820 17760
rect 480900 18348 480952 18400
rect 352684 17624 352736 17676
rect 480816 18264 480868 18316
rect 353392 17452 353444 17504
rect 12613 16017 12665 16069
rect 31212 16020 31264 16072
rect 12725 15933 12777 15985
rect 31296 15936 31348 15988
rect 12837 15849 12889 15901
rect 31380 15852 31432 15904
rect 12949 15765 13001 15817
rect 31464 15768 31516 15820
rect 13061 15681 13113 15733
rect 31548 15684 31600 15736
rect 367945 15732 368062 15849
rect 13173 15597 13225 15649
rect 31632 15600 31684 15652
rect 13960 15509 14012 15561
rect 31716 15516 31768 15568
rect 14072 15425 14124 15477
rect 31800 15432 31852 15484
rect 14184 15341 14236 15393
rect 31884 15348 31936 15400
rect 14296 15257 14348 15309
rect 31968 15264 32020 15316
rect 14408 15173 14460 15225
rect 32052 15180 32104 15232
rect 14520 15089 14572 15141
rect 32136 15096 32188 15148
rect 14632 15005 14684 15057
rect 32220 15012 32272 15064
rect 14744 14921 14796 14973
rect 32304 14928 32356 14980
rect 14856 14837 14908 14889
rect 32388 14844 32440 14896
rect 14968 14753 15020 14805
rect 32472 14760 32524 14812
rect 15079 14669 15131 14721
rect 32556 14676 32608 14728
rect 15190 14585 15242 14637
rect 32640 14592 32692 14644
rect 15301 14501 15353 14553
rect 32724 14508 32776 14560
rect 15412 14417 15464 14469
rect 32808 14424 32860 14476
rect 15523 14333 15575 14385
rect 32892 14340 32944 14392
rect 15634 14249 15686 14301
rect 32976 14256 33028 14308
rect 15745 14165 15797 14217
rect 33060 14172 33112 14224
rect 15856 14081 15908 14133
rect 33144 14088 33196 14140
rect 16204 13998 16256 14050
rect 33228 14004 33280 14056
rect 16315 13914 16367 13966
rect 33312 13920 33364 13972
rect 16426 13830 16478 13882
rect 33396 13836 33448 13888
rect 16537 13746 16589 13798
rect 33480 13752 33532 13804
rect 16648 13662 16700 13714
rect 33564 13668 33616 13720
rect 16753 13586 16805 13638
rect 33648 13584 33700 13636
rect 18884 13504 18936 13556
rect 33732 13500 33784 13552
rect 363194 13493 363246 13545
rect 18329 13414 18381 13466
rect 33816 13416 33868 13468
rect 18440 13330 18492 13382
rect 33900 13332 33952 13384
rect 18551 13246 18603 13298
rect 33984 13248 34036 13300
rect 18662 13162 18714 13214
rect 34068 13164 34120 13216
rect 18773 13078 18825 13130
rect 34152 13080 34204 13132
rect 28516 12918 28568 12970
rect 81830 12914 81882 12966
rect 28628 12834 28680 12886
rect 81914 12830 81966 12882
rect 28740 12750 28792 12802
rect 81998 12746 82050 12798
rect 28852 12665 28904 12717
rect 82082 12662 82134 12714
rect 28964 12582 29016 12634
rect 82166 12578 82218 12630
rect 29076 12498 29128 12550
rect 82250 12494 82302 12546
rect 29188 12413 29240 12465
rect 82334 12410 82386 12462
rect 29300 12329 29352 12381
rect 82418 12326 82470 12378
rect 28404 12245 28456 12297
rect 82502 12242 82554 12294
rect 28292 12161 28344 12213
rect 82586 12158 82638 12210
rect 28180 12078 28232 12130
rect 82670 12074 82722 12126
rect 28068 11993 28120 12045
rect 82754 11990 82806 12042
rect 27956 11910 28008 11962
rect 82838 11906 82890 11958
rect 27844 11828 27896 11880
rect 82922 11822 82974 11874
rect 363280 11863 363332 11915
rect 27732 11741 27784 11793
rect 83006 11738 83058 11790
rect 27620 11658 27672 11710
rect 83090 11654 83142 11706
rect 29857 11578 29909 11630
rect 80949 11578 81001 11630
rect 30646 11494 30698 11546
rect 81033 11494 81085 11546
rect 30532 11410 30584 11462
rect 81117 11410 81169 11462
rect 30308 11326 30360 11378
rect 81201 11326 81253 11378
rect 30417 11242 30469 11294
rect 81285 11242 81337 11294
rect 30978 11158 31030 11210
rect 81369 11158 81421 11210
rect 30869 11074 30921 11126
rect 81453 11074 81505 11126
rect 31430 10990 31482 11042
rect 81537 10990 81589 11042
rect 30756 10906 30808 10958
rect 81621 10906 81673 10958
rect 92028 10930 92080 10982
rect 93466 10930 93518 10982
rect 95094 10930 95146 10982
rect 96722 10930 96774 10982
rect 98350 10930 98402 10982
rect 99978 10930 100030 10982
rect 101606 10930 101658 10982
rect 103234 10930 103286 10982
rect 104862 10930 104914 10982
rect 110109 10928 110167 10986
rect 111737 10928 111795 10986
rect 113365 10928 113423 10986
rect 114993 10928 115051 10986
rect 116621 10928 116679 10986
rect 118249 10928 118307 10986
rect 119877 10928 119935 10986
rect 121505 10928 121563 10986
rect 31202 10822 31254 10874
rect 81705 10822 81757 10874
rect 23028 10746 23080 10798
rect 23140 10655 23192 10707
rect 23252 10574 23304 10626
rect 23364 10493 23416 10545
rect 23476 10404 23528 10456
rect 23588 10321 23640 10373
rect 121505 10319 121563 10377
rect 23700 10236 23752 10288
rect 119877 10229 119935 10287
rect 23812 10152 23864 10204
rect 118248 10155 118300 10207
rect 23924 10072 23976 10124
rect 116620 10067 116672 10119
rect 24036 9989 24088 10041
rect 114992 9988 115044 10040
rect 24148 9904 24200 9956
rect 113364 9904 113416 9956
rect 24260 9818 24312 9870
rect 111736 9818 111788 9870
rect 24372 9735 24424 9787
rect 110108 9733 110160 9785
rect 24484 9650 24536 9702
rect 92028 9646 92080 9698
rect 24596 9568 24648 9620
rect 24708 9480 24760 9532
rect 24820 9399 24872 9451
rect 24932 9314 24984 9366
rect 25044 9230 25096 9282
rect 93466 9226 93518 9278
rect 25156 9146 25208 9198
rect 95094 9143 95146 9195
rect 25268 9061 25320 9113
rect 96722 9055 96774 9107
rect 530536 21213 530588 21265
rect 541027 21213 541079 21265
rect 530620 21129 530672 21181
rect 541111 21129 541163 21181
rect 530704 21045 530756 21097
rect 541195 21045 541247 21097
rect 530788 20961 530840 21013
rect 541279 20961 541331 21013
rect 530872 20877 530924 20929
rect 541363 20877 541415 20929
rect 530956 20793 531008 20845
rect 541447 20793 541499 20845
rect 531040 20709 531092 20761
rect 541531 20709 541583 20761
rect 531124 20625 531176 20677
rect 541615 20625 541667 20677
rect 531208 20541 531260 20593
rect 541699 20541 541751 20593
rect 531292 20457 531344 20509
rect 541783 20457 541835 20509
rect 531376 20373 531428 20425
rect 541867 20373 541919 20425
rect 531460 20289 531512 20341
rect 541951 20289 542003 20341
rect 531544 20205 531596 20257
rect 542035 20205 542087 20257
rect 531628 20121 531680 20173
rect 542119 20121 542171 20173
rect 531712 20037 531764 20089
rect 542203 20037 542255 20089
rect 531796 19953 531848 20005
rect 542287 19953 542339 20005
rect 531880 19869 531932 19921
rect 542371 19869 542423 19921
rect 531964 19785 532016 19837
rect 542455 19785 542507 19837
rect 532048 19701 532100 19753
rect 542539 19701 542591 19753
rect 532132 19617 532184 19669
rect 542623 19617 542675 19669
rect 532216 19533 532268 19585
rect 542707 19533 542759 19585
rect 532300 19449 532352 19501
rect 542791 19449 542843 19501
rect 532384 19365 532436 19417
rect 542875 19365 542927 19417
rect 532468 19281 532520 19333
rect 542959 19281 543011 19333
rect 532552 19197 532604 19249
rect 543043 19197 543095 19249
rect 532636 19113 532688 19165
rect 543127 19113 543179 19165
rect 532720 19029 532772 19081
rect 543211 19029 543263 19081
rect 532804 18945 532856 18997
rect 543295 18945 543347 18997
rect 532888 18861 532940 18913
rect 543379 18861 543431 18913
rect 532972 18777 533024 18829
rect 543463 18777 543515 18829
rect 533056 18693 533108 18745
rect 543547 18693 543599 18745
rect 533140 18609 533192 18661
rect 543631 18609 543683 18661
rect 533224 18525 533276 18577
rect 543715 18525 543767 18577
rect 533308 18441 533360 18493
rect 543799 18441 543851 18493
rect 530258 18315 530310 18367
rect 538148 18314 538200 18366
rect 530174 18231 530226 18283
rect 538036 18230 538088 18282
rect 530090 18147 530142 18199
rect 537924 18146 537976 18198
rect 530006 18063 530058 18115
rect 537812 18062 537864 18114
rect 529922 17979 529974 18031
rect 537700 17978 537752 18030
rect 529838 17895 529890 17947
rect 537588 17894 537640 17946
rect 529754 17811 529806 17863
rect 537476 17810 537528 17862
rect 529670 17727 529722 17779
rect 537364 17726 537416 17778
rect 529586 17643 529638 17695
rect 537252 17642 537304 17694
rect 529502 17559 529554 17611
rect 537140 17558 537192 17610
rect 529418 17475 529470 17527
rect 537028 17474 537080 17526
rect 529334 17391 529386 17443
rect 536916 17390 536968 17442
rect 490687 9730 490755 9798
rect 536692 17080 536744 17132
rect 536580 16996 536632 17048
rect 536468 16912 536520 16964
rect 536356 16828 536408 16880
rect 536244 16744 536296 16796
rect 536132 16660 536184 16712
rect 536020 16576 536072 16628
rect 535908 16492 535960 16544
rect 535796 16408 535848 16460
rect 521032 14176 521084 14228
rect 520948 14052 521000 14104
rect 520860 13936 520912 13988
rect 520776 13816 520828 13868
rect 535684 16324 535736 16376
rect 535572 16240 535624 16292
rect 535460 16156 535512 16208
rect 535348 16072 535400 16124
rect 524418 15786 524470 15838
rect 553380 15790 553432 15842
rect 524334 15702 524386 15754
rect 553268 15704 553320 15756
rect 524250 15618 524302 15670
rect 552932 15622 552984 15674
rect 524166 15534 524218 15586
rect 552484 15540 552536 15592
rect 524082 15450 524134 15502
rect 552148 15452 552200 15504
rect 523998 15366 524050 15418
rect 551140 15370 551192 15422
rect 523914 15282 523966 15334
rect 551028 15288 551080 15340
rect 523830 15198 523882 15250
rect 550692 15202 550744 15254
rect 523746 15114 523798 15166
rect 550132 15118 550184 15170
rect 523662 15030 523714 15082
rect 549796 15040 549848 15092
rect 523578 14946 523630 14998
rect 545428 14954 545480 15006
rect 523494 14862 523546 14914
rect 544644 14870 544696 14922
rect 523410 14778 523462 14830
rect 543972 14780 544024 14832
rect 523326 14694 523378 14746
rect 543188 14700 543240 14752
rect 529042 14392 529094 14444
rect 528958 14318 529010 14370
rect 528874 14244 528926 14296
rect 528790 14170 528842 14222
rect 528706 14096 528758 14148
rect 528622 14022 528674 14074
rect 528538 13948 528590 14000
rect 528454 13874 528506 13926
rect 528370 13800 528422 13852
rect 528286 13726 528338 13778
rect 528202 13652 528254 13704
rect 528118 13578 528170 13630
rect 528034 13504 528086 13556
rect 527950 13430 528002 13482
rect 527866 13356 527918 13408
rect 527782 13282 527834 13334
rect 527698 13208 527750 13260
rect 527614 13134 527666 13186
rect 527530 13060 527582 13112
rect 527446 12986 527498 13038
rect 527362 12912 527414 12964
rect 527278 12838 527330 12890
rect 527194 12764 527246 12816
rect 527110 12690 527162 12742
rect 527026 12616 527078 12668
rect 526942 12542 526994 12594
rect 526858 12468 526910 12520
rect 526774 12394 526826 12446
rect 526690 12320 526742 12372
rect 526606 12246 526658 12298
rect 526522 12172 526574 12224
rect 526438 12098 526490 12150
rect 526354 12024 526406 12076
rect 526270 11950 526322 12002
rect 526186 11876 526238 11928
rect 526102 11802 526154 11854
rect 526018 11728 526070 11780
rect 525934 11654 525986 11706
rect 520698 11584 520750 11636
rect 525850 11580 525902 11632
rect 520612 11464 520664 11516
rect 525766 11506 525818 11558
rect 525682 11432 525734 11484
rect 520526 11344 520578 11396
rect 525598 11358 525650 11410
rect 525514 11284 525566 11336
rect 520442 11224 520494 11276
rect 525430 11210 525482 11262
rect 525346 11136 525398 11188
rect 525262 11062 525314 11114
rect 525178 10988 525230 11040
rect 525094 10914 525146 10966
rect 525010 10840 525062 10892
rect 524926 10766 524978 10818
rect 524842 10692 524894 10744
rect 524758 10618 524810 10670
rect 524674 10544 524726 10596
rect 534788 10328 534840 10380
rect 535236 10243 535288 10295
rect 535124 10159 535176 10211
rect 535012 10075 535064 10127
rect 534900 9989 534952 10041
rect 522955 9878 523007 9930
rect 539940 9880 539992 9932
rect 522871 9794 522923 9846
rect 539828 9796 539880 9848
rect 522787 9710 522839 9762
rect 539716 9712 539768 9764
rect 522703 9626 522755 9678
rect 539604 9628 539656 9680
rect 522619 9542 522671 9594
rect 539492 9544 539544 9596
rect 522535 9458 522587 9510
rect 539380 9460 539432 9512
rect 522451 9374 522503 9426
rect 539268 9376 539320 9428
rect 522367 9290 522419 9342
rect 539156 9292 539208 9344
rect 522283 9206 522335 9258
rect 539044 9208 539096 9260
rect 522199 9122 522251 9174
rect 538932 9124 538984 9176
rect 522115 9038 522167 9090
rect 538820 9040 538872 9092
rect 25380 8979 25432 9031
rect 98350 8971 98402 9023
rect 522031 8954 522083 9006
rect 538708 8956 538760 9008
rect 25492 8895 25544 8947
rect 99978 8887 100030 8939
rect 521947 8870 521999 8922
rect 538596 8872 538648 8924
rect 25604 8811 25656 8863
rect 101606 8803 101658 8855
rect 521863 8786 521915 8838
rect 538484 8788 538536 8840
rect 25716 8727 25768 8779
rect 103234 8719 103286 8771
rect 521779 8702 521831 8754
rect 538372 8704 538424 8756
rect 25828 8644 25880 8696
rect 104862 8641 104914 8693
rect 521695 8618 521747 8670
rect 538260 8619 538312 8671
rect 484692 8480 484744 8532
rect 542622 8480 542674 8532
rect 484608 8396 484660 8448
rect 542510 8396 542562 8448
rect 484524 8312 484576 8364
rect 542398 8312 542450 8364
rect 484440 8228 484492 8280
rect 542286 8228 542338 8280
rect 484356 8144 484408 8196
rect 542174 8144 542226 8196
rect 484272 8060 484324 8112
rect 542062 8060 542114 8112
rect 484188 7976 484240 8028
rect 541950 7976 542002 8028
rect 484104 7892 484156 7944
rect 541838 7892 541890 7944
rect 25940 7820 25992 7872
rect 233042 7814 233094 7866
rect 484020 7808 484072 7860
rect 541726 7808 541778 7860
rect 26052 7736 26104 7788
rect 173952 7730 174004 7782
rect 483936 7724 483988 7776
rect 541618 7724 541670 7776
rect 483852 7640 483904 7692
rect 541510 7640 541562 7692
rect 483768 7556 483820 7608
rect 541402 7556 541454 7608
rect 483684 7472 483736 7524
rect 541290 7472 541342 7524
rect 483600 7388 483652 7440
rect 541178 7388 541230 7440
rect 483516 7304 483568 7356
rect 541066 7304 541118 7356
rect 483432 7220 483484 7272
rect 540954 7220 541006 7272
rect 483348 7136 483400 7188
rect 540840 7136 540892 7188
rect 483264 7052 483316 7104
rect 540726 7052 540778 7104
rect 483180 6968 483232 7020
rect 540612 6968 540664 7020
rect 483096 6884 483148 6936
rect 540498 6884 540550 6936
rect 483012 6800 483064 6852
rect 540384 6800 540436 6852
rect 17316 6726 17368 6778
rect 34596 6726 34648 6778
rect 17652 6641 17704 6693
rect 34680 6642 34732 6694
rect 17764 6556 17816 6608
rect 34764 6558 34816 6610
rect 18100 6472 18152 6524
rect 34848 6474 34900 6526
rect 18212 6388 18264 6440
rect 34932 6390 34984 6442
rect 19444 6304 19496 6356
rect 35016 6306 35068 6358
rect 19780 6222 19832 6274
rect 35100 6222 35152 6274
rect 19892 6133 19944 6185
rect 35184 6138 35236 6190
rect 20228 6050 20280 6102
rect 35268 6054 35320 6106
rect 20340 5970 20392 6022
rect 35352 5970 35404 6022
rect 20900 5887 20952 5939
rect 35436 5886 35488 5938
rect 21124 5802 21176 5854
rect 35520 5802 35572 5854
rect 13284 5565 13336 5617
rect 13396 5480 13448 5532
rect 13508 5396 13560 5448
rect 13620 5312 13672 5364
rect 13732 5228 13784 5280
rect 13844 5145 13896 5197
rect 15972 5060 16024 5112
rect 16084 4978 16136 5030
rect 16868 4894 16920 4946
rect 16980 4808 17032 4860
rect 17092 4723 17144 4775
rect 17204 4642 17256 4694
rect 17428 4557 17480 4609
rect 17540 4473 17592 4525
rect 17876 4305 17928 4357
rect 17988 4220 18040 4272
rect 18996 4136 19048 4188
rect 19108 4053 19160 4105
rect 19220 3969 19272 4021
rect 19332 3885 19384 3937
rect 19556 3802 19608 3854
rect 19668 3717 19720 3769
rect 20004 3632 20056 3684
rect 20116 3548 20168 3600
rect 21012 3464 21064 3516
rect 21236 3380 21288 3432
rect 21348 3296 21400 3348
rect 21460 3212 21512 3264
rect 29412 3129 29464 3181
rect 29524 3045 29576 3097
rect 29636 2960 29688 3012
rect 29748 2876 29800 2928
rect 21572 2719 21624 2771
rect 83290 2717 83342 2769
rect 21684 2635 21736 2687
rect 83374 2633 83426 2685
rect 21796 2551 21848 2603
rect 83458 2549 83510 2601
rect 21908 2467 21960 2519
rect 83542 2465 83594 2517
rect 31561 2337 31835 2411
rect 83665 2337 83739 2611
rect 290025 5280 290077 5332
rect 543300 5285 543352 5337
rect 289941 5196 289993 5248
rect 544084 5199 544136 5251
rect 289857 5112 289909 5164
rect 544756 5115 544808 5167
rect 286725 5010 286777 5062
rect 289773 5028 289825 5080
rect 545540 5032 545592 5084
rect 286809 4926 286861 4978
rect 289689 4944 289741 4996
rect 549348 4949 549400 5001
rect 286893 4842 286945 4894
rect 289605 4860 289657 4912
rect 549460 4865 549512 4917
rect 286977 4758 287029 4810
rect 289521 4776 289573 4828
rect 549572 4782 549624 4834
rect 248005 4674 248057 4726
rect 289437 4692 289489 4744
rect 549684 4697 549736 4749
rect 248089 4590 248141 4642
rect 289353 4608 289405 4660
rect 549908 4614 549960 4666
rect 248173 4506 248225 4558
rect 289269 4524 289321 4576
rect 550020 4528 550072 4580
rect 248257 4422 248309 4474
rect 289185 4440 289237 4492
rect 550804 4445 550856 4497
rect 287061 4338 287113 4390
rect 289101 4356 289153 4408
rect 550916 4362 550968 4414
rect 287145 4254 287197 4306
rect 289017 4272 289069 4324
rect 551700 4275 551752 4327
rect 287229 4170 287281 4222
rect 288933 4188 288985 4240
rect 551812 4192 551864 4244
rect 287313 4086 287365 4138
rect 288849 4104 288901 4156
rect 551924 4108 551976 4160
rect 248677 4002 248729 4054
rect 288765 4020 288817 4072
rect 552036 4024 552088 4076
rect 248761 3918 248813 3970
rect 288681 3936 288733 3988
rect 552260 3941 552312 3993
rect 288597 3852 288649 3904
rect 552372 3856 552424 3908
rect 248929 3750 248981 3802
rect 288513 3768 288565 3820
rect 553044 3772 553096 3824
rect 249013 3666 249065 3718
rect 288429 3684 288481 3736
rect 553156 3690 553208 3742
rect 287397 3582 287449 3634
rect 288345 3600 288397 3652
rect 553940 3604 553992 3656
rect 287481 3498 287533 3550
rect 288261 3516 288313 3568
rect 554052 3520 554104 3572
rect 287565 3414 287617 3466
rect 288177 3432 288229 3484
rect 554164 3436 554216 3488
rect 287649 3330 287701 3382
rect 288093 3348 288145 3400
rect 554276 3352 554328 3404
rect 249433 3246 249485 3298
rect 288009 3264 288061 3316
rect 554388 3269 554440 3321
rect 249517 3162 249569 3214
rect 287925 3180 287977 3232
rect 554500 3185 554552 3237
rect 249601 3078 249653 3130
rect 287841 3096 287893 3148
rect 554948 3102 555000 3154
rect 249685 2994 249737 3046
rect 287757 3012 287809 3064
rect 555060 3016 555112 3068
rect 249769 2911 249821 2963
rect 363196 2882 363248 2934
rect 249853 2827 249905 2879
rect 490687 2870 490755 2938
rect 534676 2885 534728 2937
rect 467249 2798 467301 2850
rect 534564 2801 534616 2853
rect 249937 2742 249989 2794
rect 467128 2714 467180 2766
rect 534452 2717 534504 2769
rect 250021 2658 250073 2710
rect 467015 2630 467067 2682
rect 534340 2633 534392 2685
rect 286389 2574 286441 2626
rect 466894 2546 466946 2598
rect 534228 2549 534280 2601
rect 286473 2491 286525 2543
rect 469841 2462 469893 2514
rect 534116 2465 534168 2517
rect 286557 2406 286609 2458
rect 469603 2378 469655 2430
rect 534004 2381 534056 2433
rect 286641 2323 286693 2375
rect 469480 2294 469532 2346
rect 533892 2297 533944 2349
rect 22244 2215 22296 2267
rect 472313 2210 472365 2262
rect 533780 2213 533832 2265
rect 22356 2131 22408 2183
rect 194593 2129 194645 2181
rect 472437 2126 472489 2178
rect 533668 2129 533720 2181
rect 22468 2047 22520 2099
rect 197076 2044 197128 2096
rect 472191 2042 472243 2094
rect 533556 2045 533608 2097
rect 22580 1963 22632 2015
rect 472073 1958 472125 2010
rect 533444 1961 533496 2013
rect 22692 1879 22744 1931
rect 135654 1877 135706 1929
rect 474907 1874 474959 1926
rect 533332 1877 533384 1929
rect 22804 1795 22856 1847
rect 138110 1792 138162 1844
rect 475028 1790 475080 1842
rect 533220 1793 533272 1845
rect 22916 1711 22968 1763
rect 189217 1709 189269 1761
rect 474785 1706 474837 1758
rect 533108 1709 533160 1761
rect 20449 1625 20501 1677
rect 273400 1626 273452 1678
rect 474664 1622 474716 1674
rect 532996 1625 533048 1677
rect 20561 1541 20613 1593
rect 273484 1542 273536 1594
rect 477498 1538 477550 1590
rect 532884 1541 532936 1593
rect 20678 1457 20730 1509
rect 273568 1458 273620 1510
rect 469722 1454 469774 1506
rect 532772 1457 532824 1509
rect 20790 1373 20842 1425
rect 273652 1374 273704 1426
rect 482804 1370 482856 1422
rect 532660 1373 532712 1425
rect 482561 1286 482613 1338
rect 532548 1289 532600 1341
rect 477614 1202 477666 1254
rect 532436 1205 532488 1257
rect 477379 1118 477431 1170
rect 532324 1121 532376 1173
rect 477258 1034 477310 1086
rect 532212 1037 532264 1089
rect 482445 950 482497 1002
rect 532100 953 532152 1005
rect 482685 866 482737 918
rect 531988 869 532040 921
rect 480091 782 480143 834
rect 531876 785 531928 837
rect 480207 698 480259 750
rect 531764 701 531816 753
rect 479966 614 480018 666
rect 531652 617 531704 669
rect 479847 530 479899 582
rect 531540 533 531592 585
rect 363277 446 363329 498
rect 531428 449 531480 501
<< metal2 >>
rect 10608 109066 10636 109071
rect 10720 108990 10748 108993
rect 10832 108917 10860 108933
rect 2420 65287 2548 96911
rect 2716 68192 2844 96821
rect 3012 65287 3140 102726
rect 3308 67712 3436 102624
rect 3604 65287 3732 102726
rect 3900 67231 4028 95978
rect 4196 65287 4324 102239
rect 4492 66701 4620 101842
rect 4788 65287 4916 102239
rect 5084 66221 5212 95691
rect 5380 65287 5508 101927
rect 5676 65691 5804 101547
rect 5972 65287 6100 101927
rect 10148 84104 10200 84110
rect 10148 84046 10200 84052
rect 9924 78194 9976 78200
rect 9924 78136 9976 78142
rect 9700 77953 9752 77959
rect 9700 77895 9752 77901
rect 2420 65223 6102 65287
rect 2420 64832 2511 65223
rect 2431 64731 2511 64832
rect 5983 64731 6102 65223
rect 2431 64677 6102 64731
rect 9252 55895 9304 55901
rect 9252 55837 9304 55843
rect 9028 49986 9080 49992
rect 9028 49928 9080 49934
rect 8804 49749 8856 49755
rect 8804 49691 8856 49697
rect 8356 41908 8408 41915
rect 8356 41850 8408 41856
rect 7908 35997 7960 36003
rect 7908 35939 7960 35945
rect 7460 27718 7512 27724
rect 7460 27660 7512 27666
rect 7236 21796 7288 21802
rect 7236 21738 7288 21744
rect 7012 21564 7064 21570
rect 7012 21506 7064 21512
rect 7024 0 7052 21506
rect 7124 21443 7176 21449
rect 7124 21385 7176 21391
rect 7136 0 7164 21385
rect 7248 0 7276 21738
rect 7348 21677 7400 21683
rect 7348 21619 7400 21625
rect 7360 0 7388 21619
rect 7472 0 7500 27660
rect 7572 27592 7624 27598
rect 7572 27534 7624 27540
rect 7584 0 7612 27534
rect 7696 27471 7724 27484
rect 7684 27465 7736 27471
rect 7684 27407 7736 27413
rect 7696 0 7724 27407
rect 7808 27348 7836 27360
rect 7796 27342 7848 27348
rect 7796 27284 7848 27290
rect 7808 0 7836 27284
rect 7920 0 7948 35939
rect 8020 35876 8072 35882
rect 8020 35818 8072 35824
rect 8032 0 8060 35818
rect 8132 35758 8184 35764
rect 8132 35700 8184 35706
rect 8144 0 8172 35700
rect 8244 35633 8296 35639
rect 8244 35575 8296 35581
rect 8256 0 8284 35575
rect 8368 0 8396 41850
rect 8468 41783 8520 41789
rect 8468 41725 8520 41731
rect 8480 0 8508 41725
rect 8580 41658 8632 41664
rect 8580 41600 8632 41606
rect 8592 0 8620 41600
rect 8692 41543 8744 41549
rect 8692 41485 8744 41491
rect 8704 0 8732 41485
rect 8816 0 8844 49691
rect 8916 49633 8968 49639
rect 8916 49575 8968 49581
rect 8928 0 8956 49575
rect 9040 0 9068 49928
rect 9140 49876 9192 49882
rect 9140 49818 9192 49824
rect 9152 0 9180 49818
rect 9264 0 9292 55837
rect 9364 55768 9416 55774
rect 9364 55710 9416 55716
rect 9376 0 9404 55710
rect 9488 55669 9516 55674
rect 9476 55663 9528 55669
rect 9476 55605 9528 55611
rect 9488 0 9516 55605
rect 9600 55551 9628 55554
rect 9589 55545 9641 55551
rect 9589 55487 9641 55493
rect 9600 0 9628 55487
rect 9712 0 9740 77895
rect 9812 77829 9864 77835
rect 9812 77771 9864 77777
rect 9824 0 9852 77771
rect 9936 0 9964 78136
rect 10036 78065 10088 78071
rect 10036 78007 10088 78013
rect 10048 0 10076 78007
rect 10160 0 10188 84046
rect 10260 83978 10312 83984
rect 10260 83920 10312 83926
rect 10272 0 10300 83920
rect 10372 83856 10424 83862
rect 10372 83798 10424 83804
rect 10384 0 10412 83798
rect 10484 83741 10536 83747
rect 10484 83683 10536 83689
rect 10496 0 10524 83683
rect 10608 0 10636 108874
rect 10944 108840 10972 108860
rect 10720 0 10748 108798
rect 11056 108766 11084 108777
rect 10832 0 10860 108725
rect 11168 108699 11196 108714
rect 10944 0 10972 108648
rect 11280 108629 11308 108638
rect 11056 0 11084 108574
rect 11392 108560 11420 108565
rect 11168 0 11196 108507
rect 11728 108477 11756 108486
rect 11280 0 11308 108437
rect 11840 108408 11868 108427
rect 11392 0 11420 108368
rect 11952 108330 11980 108357
rect 11728 0 11756 108285
rect 12064 108264 12092 108281
rect 11840 0 11868 108216
rect 12176 108193 12204 108204
rect 11952 0 11980 108138
rect 12288 108119 12316 108138
rect 12064 0 12092 108072
rect 12400 108042 12428 108072
rect 12176 0 12204 108001
rect 12512 107968 12540 107985
rect 12288 0 12316 107927
rect 12400 0 12428 107850
rect 12512 0 12540 107776
rect 13454 96131 13670 110738
rect 13954 102008 14170 111976
rect 14354 107874 14570 112620
rect 43556 107861 43772 109514
rect 44156 101982 44372 110122
rect 44656 96113 44872 111334
rect 48434 104470 48440 104550
rect 48520 104524 48528 104550
rect 48520 104470 48633 104524
rect 48505 104468 48633 104470
rect 45408 102600 45444 102604
rect 45400 102594 45452 102600
rect 45400 102536 45452 102542
rect 45324 102516 45360 102529
rect 45316 102510 45368 102516
rect 45316 102452 45368 102458
rect 45240 102432 45276 102449
rect 45232 102426 45284 102432
rect 45232 102368 45284 102374
rect 45156 102349 45192 102366
rect 45148 102343 45200 102349
rect 45148 102285 45200 102291
rect 45072 102264 45108 102270
rect 45064 102258 45116 102264
rect 45064 102200 45116 102206
rect 44988 102179 45024 102197
rect 44980 102173 45032 102179
rect 44980 102115 45032 102121
rect 27212 89510 28184 90276
rect 44988 89308 45024 102115
rect 31220 89272 45024 89308
rect 28901 77381 28929 77390
rect 28889 77375 28941 77381
rect 28889 77317 28941 77323
rect 19170 76684 20140 77182
rect 23760 76980 24730 77168
rect 27214 76260 28184 77124
rect 27368 61276 28340 61608
rect 19326 48816 20296 48958
rect 23916 48794 24886 48954
rect 27370 48428 28340 48934
rect 27368 47314 28340 47646
rect 19326 34608 20296 34952
rect 23916 34852 24886 34976
rect 27370 34146 28340 34944
rect 19326 33076 20298 33506
rect 23916 33094 24888 33354
rect 27368 33076 28340 33874
rect 16160 20760 16482 20798
rect 24192 20792 24514 20798
rect 19588 20776 19910 20782
rect 15874 18216 16844 20760
rect 19326 20006 20296 20776
rect 23916 18810 24886 20792
rect 27680 20784 28002 20812
rect 27370 19412 28340 20784
rect 28901 17057 28929 77317
rect 28985 77297 29013 77306
rect 28973 77291 29025 77297
rect 28973 77233 29025 77239
rect 26288 17029 28929 17057
rect 12624 16075 12652 16082
rect 12613 16069 12665 16075
rect 12613 16011 12665 16017
rect 12624 0 12652 16011
rect 12725 15985 12777 15991
rect 12725 15927 12777 15933
rect 12736 0 12764 15927
rect 12837 15901 12889 15907
rect 12837 15843 12889 15849
rect 12848 0 12876 15843
rect 12949 15817 13001 15823
rect 12949 15759 13001 15765
rect 12960 0 12988 15759
rect 13061 15733 13113 15739
rect 13061 15675 13113 15681
rect 13072 0 13100 15675
rect 13184 15655 13212 15660
rect 13173 15649 13225 15655
rect 13173 15591 13225 15597
rect 13184 0 13212 15591
rect 13968 15567 13996 15574
rect 13960 15561 14012 15567
rect 13960 15503 14012 15509
rect 13284 5617 13336 5623
rect 13284 5559 13336 5565
rect 13296 0 13324 5559
rect 13396 5532 13448 5538
rect 13396 5474 13448 5480
rect 13408 0 13436 5474
rect 13508 5448 13560 5454
rect 13508 5390 13560 5396
rect 13520 0 13548 5390
rect 13620 5364 13672 5370
rect 13620 5306 13672 5312
rect 13632 0 13660 5306
rect 13732 5280 13784 5286
rect 13732 5222 13784 5228
rect 13744 0 13772 5222
rect 13844 5197 13896 5203
rect 13844 5139 13896 5145
rect 13856 0 13884 5139
rect 13968 0 13996 15503
rect 14072 15477 14124 15483
rect 14072 15419 14124 15425
rect 14080 0 14108 15419
rect 14192 15399 14220 15406
rect 14184 15393 14236 15399
rect 14184 15335 14236 15341
rect 14192 0 14220 15335
rect 14304 15315 14332 15318
rect 14296 15309 14348 15315
rect 14296 15251 14348 15257
rect 14304 0 14332 15251
rect 14408 15225 14460 15231
rect 14408 15167 14460 15173
rect 14416 0 14444 15167
rect 14528 15147 14556 15148
rect 14520 15141 14572 15147
rect 14520 15083 14572 15089
rect 14528 0 14556 15083
rect 14640 15063 14668 15068
rect 14632 15057 14684 15063
rect 14632 14999 14684 15005
rect 14640 0 14668 14999
rect 14744 14973 14796 14979
rect 14744 14915 14796 14921
rect 14752 0 14780 14915
rect 14864 14895 14892 14902
rect 14856 14889 14908 14895
rect 14856 14831 14908 14837
rect 14864 0 14892 14831
rect 14968 14805 15020 14811
rect 14968 14747 15020 14753
rect 14976 0 15004 14747
rect 15079 14721 15131 14727
rect 15079 14663 15131 14669
rect 15088 0 15116 14663
rect 15190 14637 15242 14643
rect 15190 14579 15242 14585
rect 15200 0 15228 14579
rect 15312 14559 15340 14564
rect 15301 14553 15353 14559
rect 15301 14495 15353 14501
rect 15312 0 15340 14495
rect 15424 14475 15452 14484
rect 15412 14469 15464 14475
rect 15412 14411 15464 14417
rect 15424 0 15452 14411
rect 15536 14391 15564 14396
rect 15523 14385 15575 14391
rect 15523 14327 15575 14333
rect 15536 0 15564 14327
rect 15648 14307 15676 14320
rect 15634 14301 15686 14307
rect 15634 14243 15686 14249
rect 15648 0 15676 14243
rect 15760 14223 15788 14226
rect 15745 14217 15797 14223
rect 15745 14159 15797 14165
rect 15760 0 15788 14159
rect 15872 14139 15900 14142
rect 15856 14133 15908 14139
rect 15856 14075 15908 14081
rect 15872 0 15900 14075
rect 16208 14056 16236 14058
rect 16204 14050 16256 14056
rect 16204 13992 16256 13998
rect 15972 5112 16024 5118
rect 15972 5054 16024 5060
rect 15984 0 16012 5054
rect 16084 5030 16136 5036
rect 16084 4972 16136 4978
rect 16096 0 16124 4972
rect 16208 0 16236 13992
rect 16315 13966 16367 13972
rect 16315 13908 16367 13914
rect 16320 0 16348 13908
rect 16426 13882 16478 13888
rect 16426 13824 16478 13830
rect 16432 0 16460 13824
rect 16537 13798 16589 13804
rect 16537 13740 16589 13746
rect 16544 0 16572 13740
rect 16656 13720 16684 13728
rect 16648 13714 16700 13720
rect 16648 13656 16700 13662
rect 16656 0 16684 13656
rect 16753 13638 16805 13644
rect 16753 13580 16805 13586
rect 16768 0 16796 13580
rect 18884 13556 18936 13562
rect 18884 13498 18936 13504
rect 18336 13472 18364 13478
rect 18329 13466 18381 13472
rect 18329 13408 18381 13414
rect 17328 6784 17356 6793
rect 17316 6778 17368 6784
rect 17316 6720 17368 6726
rect 16868 4946 16920 4952
rect 16868 4888 16920 4894
rect 16880 0 16908 4888
rect 16980 4860 17032 4866
rect 16980 4802 17032 4808
rect 16992 0 17020 4802
rect 17092 4775 17144 4781
rect 17092 4717 17144 4723
rect 17104 0 17132 4717
rect 17204 4694 17256 4700
rect 17204 4636 17256 4642
rect 17216 0 17244 4636
rect 17328 0 17356 6720
rect 17664 6699 17692 6700
rect 17652 6693 17704 6699
rect 17652 6635 17704 6641
rect 17428 4609 17480 4615
rect 17428 4551 17480 4557
rect 17440 0 17468 4551
rect 17540 4525 17592 4531
rect 17540 4467 17592 4473
rect 17552 0 17580 4467
rect 17664 0 17692 6635
rect 17776 6614 17804 6628
rect 17764 6608 17816 6614
rect 17764 6550 17816 6556
rect 17776 0 17804 6550
rect 18112 6530 18140 6535
rect 18100 6524 18152 6530
rect 18100 6466 18152 6472
rect 17876 4357 17928 4363
rect 17876 4299 17928 4305
rect 17888 0 17916 4299
rect 17988 4272 18040 4278
rect 17988 4214 18040 4220
rect 18000 0 18028 4214
rect 18112 0 18140 6466
rect 18224 6446 18252 6463
rect 18212 6440 18264 6446
rect 18212 6382 18264 6388
rect 18224 0 18252 6382
rect 18336 0 18364 13408
rect 18448 13388 18476 13398
rect 18440 13382 18492 13388
rect 18440 13324 18492 13330
rect 18448 0 18476 13324
rect 18551 13298 18603 13304
rect 18551 13240 18603 13246
rect 18560 0 18588 13240
rect 18672 13220 18700 13230
rect 18662 13214 18714 13220
rect 18662 13156 18714 13162
rect 18672 0 18700 13156
rect 18784 13136 18812 13142
rect 18773 13130 18825 13136
rect 18773 13072 18825 13078
rect 18784 0 18812 13072
rect 18896 0 18924 13498
rect 23040 10804 23068 10807
rect 23028 10798 23080 10804
rect 23028 10740 23080 10746
rect 19456 6362 19484 6367
rect 19444 6356 19496 6362
rect 19444 6298 19496 6304
rect 18996 4188 19048 4194
rect 18996 4130 19048 4136
rect 19008 0 19036 4130
rect 19108 4105 19160 4111
rect 19108 4047 19160 4053
rect 19120 0 19148 4047
rect 19232 4027 19260 4030
rect 19220 4021 19272 4027
rect 19220 3963 19272 3969
rect 19232 0 19260 3963
rect 19332 3937 19384 3943
rect 19332 3879 19384 3885
rect 19344 0 19372 3879
rect 19456 0 19484 6298
rect 19792 6280 19820 6288
rect 19780 6274 19832 6280
rect 19780 6216 19832 6222
rect 19556 3854 19608 3860
rect 19556 3796 19608 3802
rect 19568 0 19596 3796
rect 19668 3769 19720 3775
rect 19668 3711 19720 3717
rect 19680 0 19708 3711
rect 19792 0 19820 6216
rect 19904 6191 19932 6198
rect 19892 6185 19944 6191
rect 19892 6127 19944 6133
rect 19904 0 19932 6127
rect 20240 6108 20268 6119
rect 20228 6102 20280 6108
rect 20228 6044 20280 6050
rect 20004 3684 20056 3690
rect 20004 3626 20056 3632
rect 20016 0 20044 3626
rect 20116 3600 20168 3606
rect 20116 3542 20168 3548
rect 20128 0 20156 3542
rect 20240 0 20268 6044
rect 20352 6028 20380 6033
rect 20340 6022 20392 6028
rect 20340 5964 20392 5970
rect 20352 0 20380 5964
rect 20912 5945 20940 5947
rect 20900 5939 20952 5945
rect 20900 5881 20952 5887
rect 20464 1683 20492 1698
rect 20449 1677 20501 1683
rect 20449 1619 20501 1625
rect 20464 0 20492 1619
rect 20576 1599 20604 1609
rect 20561 1593 20613 1599
rect 20561 1535 20613 1541
rect 20576 0 20604 1535
rect 20688 1515 20716 1520
rect 20678 1509 20730 1515
rect 20678 1451 20730 1457
rect 20688 0 20716 1451
rect 20800 1431 20828 1438
rect 20790 1425 20842 1431
rect 20790 1367 20842 1373
rect 20800 0 20828 1367
rect 20912 0 20940 5881
rect 21136 5860 21164 5865
rect 21124 5854 21176 5860
rect 21124 5796 21176 5802
rect 21012 3516 21064 3522
rect 21012 3458 21064 3464
rect 21024 0 21052 3458
rect 21136 0 21164 5796
rect 21236 3432 21288 3438
rect 21236 3374 21288 3380
rect 21248 0 21276 3374
rect 21348 3348 21400 3354
rect 21348 3290 21400 3296
rect 21360 0 21388 3290
rect 21472 3270 21500 3285
rect 21460 3264 21512 3270
rect 21460 3206 21512 3212
rect 21472 0 21500 3206
rect 21584 2777 21612 2791
rect 21572 2771 21624 2777
rect 21572 2713 21624 2719
rect 21584 0 21612 2713
rect 21696 2693 21724 2707
rect 21684 2687 21736 2693
rect 21684 2629 21736 2635
rect 21696 0 21724 2629
rect 21808 2609 21836 2623
rect 21796 2603 21848 2609
rect 21796 2545 21848 2551
rect 21808 0 21836 2545
rect 21920 2525 21948 2539
rect 21908 2519 21960 2525
rect 21908 2461 21960 2467
rect 21920 0 21948 2461
rect 22256 2273 22284 2287
rect 22244 2267 22296 2273
rect 22244 2209 22296 2215
rect 22032 0 22060 1067
rect 22144 0 22172 724
rect 22256 0 22284 2209
rect 22368 2189 22396 2203
rect 22356 2183 22408 2189
rect 22356 2125 22408 2131
rect 22368 0 22396 2125
rect 22480 2105 22508 2119
rect 22468 2099 22520 2105
rect 22468 2041 22520 2047
rect 22480 0 22508 2041
rect 22592 2021 22620 2035
rect 22580 2015 22632 2021
rect 22580 1957 22632 1963
rect 22592 0 22620 1957
rect 22704 1937 22732 1951
rect 22692 1931 22744 1937
rect 22692 1873 22744 1879
rect 22704 0 22732 1873
rect 22816 1853 22844 1867
rect 22804 1847 22856 1853
rect 22804 1789 22856 1795
rect 22816 0 22844 1789
rect 22928 1769 22956 1783
rect 22916 1763 22968 1769
rect 22916 1705 22968 1711
rect 22928 0 22956 1705
rect 23040 0 23068 10740
rect 23152 10713 23180 10723
rect 23140 10707 23192 10713
rect 23140 10649 23192 10655
rect 23152 0 23180 10649
rect 23264 10632 23292 10639
rect 23252 10626 23304 10632
rect 23252 10568 23304 10574
rect 23264 0 23292 10568
rect 23376 10551 23404 10555
rect 23364 10545 23416 10551
rect 23364 10487 23416 10493
rect 23376 0 23404 10487
rect 23488 10462 23516 10471
rect 23476 10456 23528 10462
rect 23476 10398 23528 10404
rect 23488 0 23516 10398
rect 23600 10379 23628 10387
rect 23588 10373 23640 10379
rect 23588 10315 23640 10321
rect 23600 0 23628 10315
rect 23712 10294 23740 10303
rect 23700 10288 23752 10294
rect 23700 10230 23752 10236
rect 23712 0 23740 10230
rect 23824 10204 23852 10219
rect 23806 10152 23812 10204
rect 23864 10152 23870 10204
rect 23824 0 23852 10152
rect 23936 10124 23964 10135
rect 23918 10072 23924 10124
rect 23976 10072 23982 10124
rect 23936 0 23964 10072
rect 24048 10047 24076 10051
rect 24036 10041 24088 10047
rect 24036 9983 24088 9989
rect 24048 0 24076 9983
rect 24160 9962 24188 9967
rect 24148 9956 24200 9962
rect 24148 9898 24200 9904
rect 24160 0 24188 9898
rect 24272 9876 24300 9883
rect 24260 9870 24312 9876
rect 24260 9812 24312 9818
rect 24272 0 24300 9812
rect 24384 9793 24412 9799
rect 24372 9787 24424 9793
rect 24372 9729 24424 9735
rect 24384 0 24412 9729
rect 24496 9708 24524 9715
rect 24484 9702 24536 9708
rect 24484 9644 24536 9650
rect 24496 0 24524 9644
rect 24608 9626 24636 9631
rect 24596 9620 24648 9626
rect 24596 9562 24648 9568
rect 24608 0 24636 9562
rect 24720 9538 24748 9547
rect 24708 9532 24760 9538
rect 24708 9474 24760 9480
rect 24720 0 24748 9474
rect 24832 9457 24860 9463
rect 24820 9451 24872 9457
rect 24820 9393 24872 9399
rect 24832 0 24860 9393
rect 24944 9372 24972 9379
rect 24932 9366 24984 9372
rect 24932 9308 24984 9314
rect 24944 0 24972 9308
rect 25056 9288 25084 9295
rect 25044 9282 25096 9288
rect 25044 9224 25096 9230
rect 25056 0 25084 9224
rect 25168 9204 25196 9211
rect 25156 9198 25208 9204
rect 25156 9140 25208 9146
rect 25168 0 25196 9140
rect 25280 9119 25308 9127
rect 25268 9113 25320 9119
rect 25268 9055 25320 9061
rect 25280 0 25308 9055
rect 25392 9037 25420 9043
rect 25380 9031 25432 9037
rect 25380 8973 25432 8979
rect 25392 0 25420 8973
rect 25504 8947 25532 8959
rect 25486 8895 25492 8947
rect 25544 8895 25550 8947
rect 25504 0 25532 8895
rect 25616 8869 25644 8875
rect 25604 8863 25656 8869
rect 25604 8805 25656 8811
rect 25616 0 25644 8805
rect 25728 8785 25756 8791
rect 25716 8779 25768 8785
rect 25716 8721 25768 8727
rect 25728 0 25756 8721
rect 25840 8702 25868 8707
rect 25828 8696 25880 8702
rect 25828 8638 25880 8644
rect 25840 0 25868 8638
rect 25952 7878 25980 7883
rect 25940 7872 25992 7878
rect 25940 7814 25992 7820
rect 25952 0 25980 7814
rect 26064 7794 26092 7799
rect 26052 7788 26104 7794
rect 26052 7730 26104 7736
rect 26064 0 26092 7730
rect 26176 0 26204 395
rect 26288 0 26316 17029
rect 28985 16973 29013 77233
rect 29069 77213 29097 77222
rect 29057 77207 29109 77213
rect 29057 77149 29109 77155
rect 26400 16945 29013 16973
rect 26400 0 26428 16945
rect 29069 16889 29097 77149
rect 29153 77129 29181 77138
rect 29141 77123 29193 77129
rect 29141 77065 29193 77071
rect 26512 16861 29097 16889
rect 26512 0 26540 16861
rect 29153 16805 29181 77065
rect 29237 77045 29265 77054
rect 29225 77039 29277 77045
rect 29225 76981 29277 76987
rect 26624 16777 29181 16805
rect 26624 0 26652 16777
rect 29237 16721 29265 76981
rect 29321 76961 29349 76970
rect 29309 76955 29361 76961
rect 29309 76897 29361 76903
rect 26736 16693 29265 16721
rect 26736 0 26764 16693
rect 29321 16637 29349 76897
rect 29405 76877 29433 76886
rect 29393 76871 29445 76877
rect 29393 76813 29445 76819
rect 26848 16609 29349 16637
rect 26848 0 26876 16609
rect 29405 16553 29433 76813
rect 29489 76793 29517 76802
rect 29477 76787 29529 76793
rect 29477 76729 29529 76735
rect 26960 16525 29433 16553
rect 26960 0 26988 16525
rect 29489 16469 29517 76729
rect 29573 76709 29601 76718
rect 29561 76703 29613 76709
rect 29561 76645 29613 76651
rect 27072 16441 29517 16469
rect 27072 0 27100 16441
rect 29573 16385 29601 76645
rect 29657 76625 29685 76634
rect 29645 76619 29697 76625
rect 29645 76561 29697 76567
rect 27184 16357 29601 16385
rect 27184 0 27212 16357
rect 29657 16301 29685 76561
rect 29741 76541 29769 76550
rect 29729 76535 29781 76541
rect 29729 76477 29781 76483
rect 27296 16273 29685 16301
rect 27296 0 27324 16273
rect 29741 16217 29769 76477
rect 29825 76457 29853 76466
rect 29813 76451 29865 76457
rect 29813 76393 29865 76399
rect 27408 16189 29769 16217
rect 27408 0 27436 16189
rect 29825 16133 29853 76393
rect 30185 57223 30213 57228
rect 30174 57217 30226 57223
rect 30174 57159 30226 57165
rect 30017 57139 30045 57149
rect 30005 57133 30057 57139
rect 30005 57075 30057 57081
rect 27520 16105 29853 16133
rect 27520 0 27548 16105
rect 30017 13643 30045 57075
rect 30101 57055 30129 57065
rect 30089 57049 30141 57055
rect 30089 56991 30141 56997
rect 30101 13768 30129 56991
rect 30185 13876 30213 57159
rect 31025 56971 31053 56980
rect 31013 56965 31065 56971
rect 31013 56907 31065 56913
rect 30857 56887 30885 56900
rect 30846 56881 30898 56887
rect 30846 56823 30898 56829
rect 30857 14772 30885 56823
rect 31025 14996 31053 56907
rect 31220 16078 31256 89272
rect 45072 89224 45108 102200
rect 31304 89188 45108 89224
rect 31212 16072 31264 16078
rect 31212 16014 31264 16020
rect 31304 15994 31340 89188
rect 45156 89140 45192 102285
rect 31388 89104 45192 89140
rect 31296 15988 31348 15994
rect 31296 15930 31348 15936
rect 31388 15910 31424 89104
rect 45240 89056 45276 102368
rect 31472 89020 45276 89056
rect 31380 15904 31432 15910
rect 31380 15846 31432 15852
rect 31388 15842 31424 15846
rect 31472 15826 31508 89020
rect 45324 88972 45360 102452
rect 31556 88936 45360 88972
rect 31464 15820 31516 15826
rect 31464 15762 31516 15768
rect 31556 15742 31592 88936
rect 45408 88888 45444 102536
rect 46920 102097 46956 102106
rect 46912 102091 46964 102097
rect 48324 102070 48330 102150
rect 48410 102148 48416 102150
rect 48410 102092 48663 102148
rect 48410 102070 48416 102092
rect 46912 102033 46964 102039
rect 46836 102013 46872 102022
rect 46828 102007 46880 102013
rect 46828 101949 46880 101955
rect 46752 101928 46788 101933
rect 46744 101922 46796 101928
rect 46744 101864 46796 101870
rect 46668 101844 46704 101850
rect 46660 101838 46712 101844
rect 46660 101780 46712 101786
rect 46584 101761 46620 101774
rect 46576 101755 46628 101761
rect 46576 101697 46628 101703
rect 46500 101678 46536 101689
rect 46492 101672 46544 101678
rect 46492 101614 46544 101620
rect 46416 96232 46452 96239
rect 46408 96226 46460 96232
rect 46408 96168 46460 96174
rect 46332 96147 46368 96156
rect 46324 96141 46376 96147
rect 46324 96083 46376 96089
rect 46248 96064 46284 96069
rect 46240 96058 46292 96064
rect 46240 96000 46292 96006
rect 46164 95978 46200 95986
rect 46156 95972 46208 95978
rect 46156 95914 46208 95920
rect 46080 95898 46116 95903
rect 46072 95892 46124 95898
rect 46072 95834 46124 95840
rect 45996 95810 46032 95824
rect 45988 95804 46040 95810
rect 45988 95746 46040 95752
rect 45912 90867 45948 90870
rect 45904 90861 45956 90867
rect 45904 90803 45956 90809
rect 45828 90786 45864 90791
rect 45820 90780 45872 90786
rect 45820 90722 45872 90728
rect 45744 90701 45780 90704
rect 45736 90695 45788 90701
rect 45736 90637 45788 90643
rect 45660 90617 45696 90622
rect 45652 90611 45704 90617
rect 45652 90553 45704 90559
rect 45576 90533 45612 90539
rect 45568 90527 45620 90533
rect 45568 90469 45620 90475
rect 45492 90449 45528 90456
rect 45484 90443 45536 90449
rect 45484 90385 45536 90391
rect 31640 88852 45444 88888
rect 31548 15736 31600 15742
rect 31548 15678 31600 15684
rect 31556 15668 31592 15678
rect 31640 15658 31676 88852
rect 45492 88804 45528 90385
rect 31724 88768 45528 88804
rect 31632 15652 31684 15658
rect 31632 15594 31684 15600
rect 31724 15574 31760 88768
rect 45576 88720 45612 90469
rect 31808 88684 45612 88720
rect 31716 15568 31768 15574
rect 31716 15510 31768 15516
rect 31808 15490 31844 88684
rect 45660 88636 45696 90553
rect 31892 88600 45696 88636
rect 31800 15484 31852 15490
rect 31800 15426 31852 15432
rect 31892 15406 31928 88600
rect 45744 88552 45780 90637
rect 31976 88516 45780 88552
rect 31884 15400 31936 15406
rect 31884 15342 31936 15348
rect 31892 15338 31928 15342
rect 31976 15322 32012 88516
rect 45828 88468 45864 90722
rect 32060 88432 45864 88468
rect 31968 15316 32020 15322
rect 31968 15258 32020 15264
rect 32060 15238 32096 88432
rect 45912 88384 45948 90803
rect 32144 88348 45948 88384
rect 32052 15232 32104 15238
rect 32052 15174 32104 15180
rect 32144 15154 32180 88348
rect 45996 88300 46032 95746
rect 32228 88264 46032 88300
rect 32136 15148 32188 15154
rect 32136 15090 32188 15096
rect 32144 15088 32180 15090
rect 32228 15070 32264 88264
rect 46080 88216 46116 95834
rect 32312 88180 46116 88216
rect 32220 15064 32272 15070
rect 32220 15006 32272 15012
rect 31025 14968 31356 14996
rect 32312 14986 32348 88180
rect 46164 88132 46200 95914
rect 32396 88096 46200 88132
rect 30857 14744 31132 14772
rect 30185 13848 30236 13876
rect 29984 13615 30045 13643
rect 30096 13736 30129 13768
rect 28528 12976 28556 12983
rect 28516 12970 28568 12976
rect 28516 12912 28568 12918
rect 28416 12303 28444 12304
rect 28404 12297 28456 12303
rect 28404 12239 28456 12245
rect 28304 12219 28332 12230
rect 28292 12213 28344 12219
rect 28292 12155 28344 12161
rect 28192 12136 28220 12143
rect 28180 12130 28232 12136
rect 28180 12072 28232 12078
rect 28080 12051 28108 12055
rect 28068 12045 28120 12051
rect 28068 11987 28120 11993
rect 27968 11968 27996 11972
rect 27956 11962 28008 11968
rect 27956 11904 28008 11910
rect 27856 11886 27884 11901
rect 27844 11880 27896 11886
rect 27844 11822 27896 11828
rect 27744 11799 27772 11810
rect 27732 11793 27784 11799
rect 27732 11735 27784 11741
rect 27632 11716 27660 11718
rect 27620 11710 27672 11716
rect 27620 11652 27672 11658
rect 27632 0 27660 11652
rect 27744 0 27772 11735
rect 27856 0 27884 11822
rect 27968 0 27996 11904
rect 28080 0 28108 11987
rect 28192 0 28220 12072
rect 28304 0 28332 12155
rect 28416 0 28444 12239
rect 28528 0 28556 12912
rect 28640 12892 28668 12898
rect 28628 12886 28680 12892
rect 28628 12828 28680 12834
rect 28640 0 28668 12828
rect 28752 12808 28780 12811
rect 28740 12802 28792 12808
rect 28740 12744 28792 12750
rect 28752 0 28780 12744
rect 28864 12723 28892 12727
rect 28852 12717 28904 12723
rect 28852 12659 28904 12665
rect 28864 0 28892 12659
rect 28976 12640 29004 12645
rect 28964 12634 29016 12640
rect 28964 12576 29016 12582
rect 28976 0 29004 12576
rect 29088 12556 29116 12559
rect 29076 12550 29128 12556
rect 29076 12492 29128 12498
rect 29088 0 29116 12492
rect 29200 12471 29228 12476
rect 29188 12465 29240 12471
rect 29188 12407 29240 12413
rect 29200 0 29228 12407
rect 29312 12387 29340 12393
rect 29300 12381 29352 12387
rect 29300 12323 29352 12329
rect 29312 0 29340 12323
rect 29872 11636 29900 11638
rect 29857 11630 29909 11636
rect 29857 11572 29909 11578
rect 29412 3181 29464 3187
rect 29412 3123 29464 3129
rect 29424 0 29452 3123
rect 29536 3103 29564 3109
rect 29524 3097 29576 3103
rect 29524 3039 29576 3045
rect 29536 0 29564 3039
rect 29648 3018 29676 3022
rect 29636 3012 29688 3018
rect 29636 2954 29688 2960
rect 29648 0 29676 2954
rect 29760 2934 29788 2937
rect 29748 2928 29800 2934
rect 29748 2870 29800 2876
rect 29760 0 29788 2870
rect 29872 0 29900 11572
rect 29984 0 30012 13615
rect 30096 0 30124 13736
rect 30208 0 30236 13848
rect 30656 11552 30684 11562
rect 30646 11546 30698 11552
rect 30646 11488 30698 11494
rect 30544 11468 30572 11475
rect 30532 11462 30584 11468
rect 30532 11404 30584 11410
rect 30320 11384 30348 11387
rect 30308 11378 30360 11384
rect 30308 11320 30360 11326
rect 30320 0 30348 11320
rect 30432 11300 30460 11311
rect 30417 11294 30469 11300
rect 30417 11236 30469 11242
rect 30432 0 30460 11236
rect 30544 0 30572 11404
rect 30656 0 30684 11488
rect 30992 11216 31020 11222
rect 30978 11210 31030 11216
rect 30978 11152 31030 11158
rect 30869 11126 30921 11132
rect 30869 11068 30921 11074
rect 30768 10964 30796 10975
rect 30756 10958 30808 10964
rect 30756 10900 30808 10906
rect 30768 0 30796 10900
rect 30880 0 30908 11068
rect 30992 0 31020 11152
rect 31104 0 31132 14744
rect 31216 10880 31244 10885
rect 31202 10874 31254 10880
rect 31202 10816 31254 10822
rect 31216 0 31244 10816
rect 31328 0 31356 14968
rect 32304 14980 32356 14986
rect 32304 14922 32356 14928
rect 32396 14902 32432 88096
rect 46248 88048 46284 96000
rect 32480 88012 46284 88048
rect 32388 14896 32440 14902
rect 32388 14838 32440 14844
rect 32480 14818 32516 88012
rect 46332 87964 46368 96083
rect 32564 87928 46368 87964
rect 32472 14812 32524 14818
rect 32472 14754 32524 14760
rect 32564 14734 32600 87928
rect 46416 87880 46452 96168
rect 32648 87844 46452 87880
rect 32556 14728 32608 14734
rect 32556 14670 32608 14676
rect 32648 14650 32684 87844
rect 46500 87796 46536 101614
rect 32732 87760 46536 87796
rect 32640 14644 32692 14650
rect 32640 14586 32692 14592
rect 32732 14566 32768 87760
rect 46584 87712 46620 101697
rect 32816 87676 46620 87712
rect 32724 14560 32776 14566
rect 32724 14502 32776 14508
rect 32816 14482 32852 87676
rect 46668 87628 46704 101780
rect 32900 87592 46704 87628
rect 32808 14476 32860 14482
rect 32808 14418 32860 14424
rect 32900 14398 32936 87592
rect 46752 87544 46788 101864
rect 32984 87508 46788 87544
rect 32892 14392 32944 14398
rect 32892 14334 32944 14340
rect 32984 14314 33020 87508
rect 46836 87460 46872 101949
rect 33068 87424 46872 87460
rect 32976 14308 33028 14314
rect 32976 14250 33028 14256
rect 33068 14230 33104 87424
rect 46920 87376 46956 102033
rect 48224 99700 48230 99780
rect 48310 99752 48316 99780
rect 48310 99700 48710 99752
rect 48298 99696 48710 99700
rect 48114 97300 48120 97380
rect 48200 97356 48213 97380
rect 48200 97300 48695 97356
rect 47416 96728 47468 96734
rect 47416 96670 47468 96676
rect 47340 96650 47376 96656
rect 47332 96644 47384 96650
rect 47332 96586 47384 96592
rect 47256 96567 47292 96571
rect 47248 96561 47300 96567
rect 47248 96503 47300 96509
rect 47172 96483 47208 96487
rect 47164 96477 47216 96483
rect 47164 96419 47216 96425
rect 47088 96397 47124 96401
rect 47080 96391 47132 96397
rect 47080 96333 47132 96339
rect 47004 96316 47040 96325
rect 46996 96310 47048 96316
rect 46996 96252 47048 96258
rect 33152 87340 46956 87376
rect 33060 14224 33112 14230
rect 33060 14166 33112 14172
rect 33152 14146 33188 87340
rect 47004 87292 47040 96252
rect 33236 87256 47040 87292
rect 33144 14140 33196 14146
rect 33144 14082 33196 14088
rect 33236 14062 33272 87256
rect 47088 87208 47124 96333
rect 33320 87172 47124 87208
rect 33228 14056 33280 14062
rect 33228 13998 33280 14004
rect 33320 13978 33356 87172
rect 47172 87124 47208 96419
rect 33404 87088 47208 87124
rect 33312 13972 33364 13978
rect 33312 13914 33364 13920
rect 33404 13894 33440 87088
rect 47256 87040 47292 96503
rect 33488 87004 47292 87040
rect 33396 13888 33448 13894
rect 33396 13830 33448 13836
rect 33488 13810 33524 87004
rect 47340 86956 47376 96586
rect 33572 86920 47376 86956
rect 33480 13804 33532 13810
rect 33480 13746 33532 13752
rect 33572 13726 33608 86920
rect 47424 86872 47460 96670
rect 48008 94900 48014 94980
rect 48094 94960 48107 94980
rect 48094 94904 48674 94960
rect 48094 94900 48107 94904
rect 88468 92894 88668 109331
rect 88876 94758 89116 111356
rect 89350 98142 89592 113219
rect 89814 102804 90082 111958
rect 91305 109069 91357 109075
rect 91305 109011 91357 109017
rect 91182 108997 91234 109003
rect 91182 108939 91234 108945
rect 91052 108925 91104 108932
rect 91052 108867 91104 108873
rect 90936 108853 90988 108859
rect 90936 108795 90988 108801
rect 90946 107729 90978 108795
rect 91069 107744 91101 108867
rect 91059 107738 91111 107744
rect 90930 107677 90936 107729
rect 90988 107677 90994 107729
rect 91192 107728 91224 108939
rect 91308 107735 91340 109011
rect 91676 108214 91930 113875
rect 102077 108934 102331 114276
rect 96965 108781 97017 108787
rect 96965 108723 97017 108729
rect 96846 108709 96898 108715
rect 96846 108651 96898 108657
rect 91298 107729 91350 107735
rect 91059 107680 91111 107686
rect 91182 107722 91234 107728
rect 96856 107717 96888 108651
rect 91298 107671 91350 107677
rect 96846 107711 96898 107717
rect 91182 107664 91234 107670
rect 96975 107705 97007 108723
rect 102077 108680 103168 108934
rect 97208 108637 97260 108643
rect 97208 108579 97260 108585
rect 97084 108565 97136 108571
rect 97084 108507 97136 108513
rect 97094 107726 97126 108507
rect 97084 107720 97136 107726
rect 96846 107653 96898 107659
rect 96965 107699 97017 107705
rect 97218 107705 97250 108579
rect 97084 107662 97136 107668
rect 97208 107699 97260 107705
rect 96965 107641 97017 107647
rect 97208 107641 97260 107647
rect 102914 106244 103168 108680
rect 102572 105990 103168 106244
rect 89814 102536 90380 102804
rect 103331 102696 103585 110056
rect 102574 102442 103585 102696
rect 89350 97900 90380 98142
rect 103883 98116 104137 114421
rect 102507 97862 104137 98116
rect 88876 94518 90366 94758
rect 104356 94704 104596 109508
rect 126088 107025 126657 110757
rect 175954 105765 176244 110571
rect 178415 105704 178703 109990
rect 228226 107276 228809 110088
rect 102588 94464 104596 94704
rect 48544 92517 48550 92569
rect 48602 92517 48668 92569
rect 47500 90360 47552 90366
rect 47500 90302 47552 90308
rect 154532 90355 156082 90383
rect 33656 86836 47460 86872
rect 33564 13720 33616 13726
rect 33564 13662 33616 13668
rect 33656 13642 33692 86836
rect 47508 86788 47544 90302
rect 47920 90274 47972 90280
rect 47920 90216 47972 90222
rect 154532 90232 154585 90355
rect 156040 90232 156082 90355
rect 47836 90190 47888 90196
rect 47836 90132 47888 90138
rect 47752 90106 47804 90112
rect 47752 90048 47804 90054
rect 47676 90028 47712 90030
rect 47668 90022 47720 90028
rect 47668 89964 47720 89970
rect 47584 89938 47636 89944
rect 47584 89880 47636 89886
rect 33740 86752 47544 86788
rect 33648 13636 33700 13642
rect 33648 13578 33700 13584
rect 33740 13558 33776 86752
rect 47592 86704 47628 89880
rect 33824 86668 47628 86704
rect 33732 13552 33784 13558
rect 33732 13494 33784 13500
rect 33824 13474 33860 86668
rect 47676 86620 47712 89964
rect 33908 86584 47712 86620
rect 33816 13468 33868 13474
rect 33816 13410 33868 13416
rect 33908 13390 33944 86584
rect 47760 86536 47796 90048
rect 33992 86500 47796 86536
rect 33900 13384 33952 13390
rect 33900 13326 33952 13332
rect 33992 13306 34028 86500
rect 47844 86452 47880 90132
rect 34076 86416 47880 86452
rect 33984 13300 34036 13306
rect 33984 13242 34036 13248
rect 34076 13222 34112 86416
rect 47928 86368 47964 90216
rect 154532 90196 156082 90232
rect 48526 90100 48532 90180
rect 48612 90164 48618 90180
rect 48612 90108 48648 90164
rect 48612 90100 48618 90108
rect 154634 88824 156048 88857
rect 154634 88696 154673 88824
rect 156003 88696 156048 88824
rect 154634 88671 156048 88696
rect 48344 87746 48673 87748
rect 48344 87694 48365 87746
rect 48417 87694 48673 87746
rect 48344 87692 48673 87694
rect 34160 86332 47964 86368
rect 34068 13216 34120 13222
rect 34068 13158 34120 13164
rect 34160 13138 34196 86332
rect 48246 85370 48673 85372
rect 48246 85318 48261 85370
rect 48313 85318 48673 85370
rect 48246 85316 48673 85318
rect 157962 83132 158140 95999
rect 196222 89886 196274 89892
rect 196222 89828 196274 89834
rect 158294 89591 158300 89643
rect 158352 89591 158358 89643
rect 48141 82910 48157 82966
rect 48213 82910 48727 82966
rect 147547 82869 158140 83132
rect 147547 81954 147810 82869
rect 147164 81522 147810 81954
rect 151632 81513 153172 81944
rect 156173 81513 157122 81944
rect 47281 81227 49082 81245
rect 47281 81226 48765 81227
rect 47281 80913 47304 81226
rect 47726 80913 48765 81226
rect 47281 80907 48765 80913
rect 49066 80907 49082 81227
rect 147166 80966 147520 81390
rect 47281 80890 49082 80907
rect 47281 79997 49082 80015
rect 47281 79996 48765 79997
rect 47281 79683 47304 79996
rect 47726 79683 48765 79996
rect 47281 79677 48765 79683
rect 49066 79677 49082 79997
rect 47281 79660 49082 79677
rect 53196 77745 53332 78528
rect 64616 77136 64816 78330
rect 74340 76386 74540 78332
rect 84034 77171 84234 78330
rect 94238 77841 94274 77846
rect 94230 77835 94282 77841
rect 94230 77777 94282 77783
rect 84034 76971 85379 77171
rect 34604 76083 34640 76088
rect 34596 76077 34648 76083
rect 34596 76019 34648 76025
rect 34152 13132 34204 13138
rect 34152 13074 34204 13080
rect 31440 11048 31468 11051
rect 31430 11042 31482 11048
rect 31430 10984 31482 10990
rect 31440 0 31468 10984
rect 34604 6784 34640 76019
rect 34688 75999 34724 76004
rect 34680 75993 34732 75999
rect 34680 75935 34732 75941
rect 34596 6778 34648 6784
rect 34596 6720 34648 6726
rect 34604 6716 34640 6720
rect 34688 6700 34724 75935
rect 34772 75915 34808 75920
rect 34764 75909 34816 75915
rect 34764 75851 34816 75857
rect 34680 6694 34732 6700
rect 34680 6636 34732 6642
rect 34688 6632 34724 6636
rect 34772 6616 34808 75851
rect 34856 75831 34892 75836
rect 34848 75825 34900 75831
rect 34848 75767 34900 75773
rect 34764 6610 34816 6616
rect 34764 6552 34816 6558
rect 34772 6548 34808 6552
rect 34856 6532 34892 75767
rect 34940 75747 34976 75752
rect 34932 75741 34984 75747
rect 34932 75683 34984 75689
rect 34848 6526 34900 6532
rect 34848 6468 34900 6474
rect 34856 6464 34892 6468
rect 34940 6448 34976 75683
rect 35024 75663 35060 75668
rect 35016 75657 35068 75663
rect 35016 75599 35068 75605
rect 34932 6442 34984 6448
rect 34932 6384 34984 6390
rect 34940 6380 34976 6384
rect 35024 6364 35060 75599
rect 35108 75579 35144 75584
rect 35100 75573 35152 75579
rect 35100 75515 35152 75521
rect 35016 6358 35068 6364
rect 35016 6300 35068 6306
rect 35024 6296 35060 6300
rect 35108 6280 35144 75515
rect 35192 75495 35228 75500
rect 35184 75489 35236 75495
rect 35184 75431 35236 75437
rect 35100 6274 35152 6280
rect 35100 6216 35152 6222
rect 35108 6212 35144 6216
rect 35192 6196 35228 75431
rect 35276 75411 35312 75416
rect 35268 75405 35320 75411
rect 35268 75347 35320 75353
rect 35184 6190 35236 6196
rect 35184 6132 35236 6138
rect 35192 6128 35228 6132
rect 35276 6112 35312 75347
rect 35360 75327 35396 75332
rect 35352 75321 35404 75327
rect 35352 75263 35404 75269
rect 35268 6106 35320 6112
rect 35268 6048 35320 6054
rect 35276 6044 35312 6048
rect 35360 6028 35396 75263
rect 35444 75243 35480 75248
rect 35436 75237 35488 75243
rect 35436 75179 35488 75185
rect 35352 6022 35404 6028
rect 35352 5964 35404 5970
rect 35360 5960 35396 5964
rect 35444 5944 35480 75179
rect 35528 75159 35564 75164
rect 35520 75153 35572 75159
rect 35520 75095 35572 75101
rect 35436 5938 35488 5944
rect 35436 5880 35488 5886
rect 35444 5876 35480 5880
rect 35528 5860 35564 75095
rect 94238 69426 94274 77777
rect 94322 77757 94358 77762
rect 94314 77751 94366 77757
rect 94314 77693 94366 77699
rect 81838 69390 94274 69426
rect 48575 56534 48639 61797
rect 52575 56595 52639 62176
rect 76404 57217 76456 57223
rect 76404 57159 76456 57165
rect 70620 57139 70648 57146
rect 70609 57133 70661 57139
rect 70609 57075 70661 57081
rect 69976 57055 70004 57063
rect 69968 57049 70020 57055
rect 69968 56991 70020 56997
rect 67370 56965 67430 56976
rect 67370 56913 67378 56965
rect 64930 56881 64986 56891
rect 64930 56829 64933 56881
rect 64985 56829 64986 56881
rect 64930 56597 64986 56829
rect 67370 56595 67430 56913
rect 69976 56636 70004 56991
rect 70620 56636 70648 57075
rect 76416 56636 76444 57159
rect 81713 49786 81749 49806
rect 81705 49777 81761 49786
rect 81705 49712 81761 49721
rect 81629 49106 81665 49129
rect 81620 49097 81676 49106
rect 81620 49032 81676 49041
rect 81545 47746 81581 47759
rect 81540 47737 81596 47746
rect 81540 47672 81596 47681
rect 81461 47066 81497 47088
rect 81451 47057 81507 47066
rect 81451 46992 81507 47001
rect 81377 45706 81413 45723
rect 81368 45697 81424 45706
rect 81368 45632 81424 45641
rect 81293 41919 81329 41936
rect 81285 41910 81341 41919
rect 81285 41845 81341 41854
rect 81209 41569 81245 41588
rect 81200 41560 81256 41569
rect 81200 41495 81256 41504
rect 81125 41261 81161 41276
rect 81116 41252 81172 41261
rect 81116 41187 81172 41196
rect 81041 39180 81077 39199
rect 81032 39171 81088 39180
rect 81032 39106 81088 39115
rect 80957 38585 80993 38604
rect 80946 38576 81002 38585
rect 80946 38511 81002 38520
rect 80957 11636 80993 38511
rect 80949 11630 81001 11636
rect 80949 11572 81001 11578
rect 80957 11568 80993 11572
rect 81041 11552 81077 39106
rect 81033 11546 81085 11552
rect 81033 11488 81085 11494
rect 81041 11484 81077 11488
rect 81125 11468 81161 41187
rect 81117 11462 81169 11468
rect 81117 11404 81169 11410
rect 81125 11400 81161 11404
rect 81209 11384 81245 41495
rect 81201 11378 81253 11384
rect 81201 11320 81253 11326
rect 81209 11316 81245 11320
rect 81293 11300 81329 41845
rect 81285 11294 81337 11300
rect 81285 11236 81337 11242
rect 81293 11232 81329 11236
rect 81377 11216 81413 45632
rect 81369 11210 81421 11216
rect 81369 11152 81421 11158
rect 81377 11148 81413 11152
rect 81461 11132 81497 46992
rect 81453 11126 81505 11132
rect 81453 11068 81505 11074
rect 81461 11064 81497 11068
rect 81545 11048 81581 47672
rect 81537 11042 81589 11048
rect 81537 10984 81589 10990
rect 81545 10980 81581 10984
rect 81629 10964 81665 49032
rect 81621 10958 81673 10964
rect 81621 10900 81673 10906
rect 81629 10896 81665 10900
rect 81713 10880 81749 49712
rect 81838 12972 81874 69390
rect 94322 69342 94358 77693
rect 94406 77673 94442 77678
rect 94398 77667 94450 77673
rect 94398 77609 94450 77615
rect 81922 69306 94358 69342
rect 81830 12966 81882 12972
rect 81830 12908 81882 12914
rect 81838 12904 81874 12908
rect 81922 12888 81958 69306
rect 94406 69258 94442 77609
rect 94490 77589 94526 77594
rect 94482 77583 94534 77589
rect 94482 77525 94534 77531
rect 82006 69222 94442 69258
rect 81914 12882 81966 12888
rect 81914 12824 81966 12830
rect 81922 12820 81958 12824
rect 82006 12804 82042 69222
rect 94490 69174 94526 77525
rect 94574 77505 94610 77510
rect 94566 77499 94618 77505
rect 94566 77441 94618 77447
rect 82090 69138 94526 69174
rect 81998 12798 82050 12804
rect 81998 12740 82050 12746
rect 82006 12736 82042 12740
rect 82090 12720 82126 69138
rect 94574 69090 94610 77441
rect 94658 77421 94694 77426
rect 94650 77415 94702 77421
rect 94650 77357 94702 77363
rect 82174 69054 94610 69090
rect 82082 12714 82134 12720
rect 82082 12656 82134 12662
rect 82090 12652 82126 12656
rect 82174 12636 82210 69054
rect 94658 69006 94694 77357
rect 94742 77337 94778 77342
rect 94734 77331 94786 77337
rect 94734 77273 94786 77279
rect 82258 68970 94694 69006
rect 82166 12630 82218 12636
rect 82166 12572 82218 12578
rect 82174 12568 82210 12572
rect 82258 12552 82294 68970
rect 94742 68922 94778 77273
rect 94826 77253 94862 77258
rect 94818 77247 94870 77253
rect 94818 77189 94870 77195
rect 82342 68886 94778 68922
rect 82250 12546 82302 12552
rect 82250 12488 82302 12494
rect 82258 12484 82294 12488
rect 82342 12468 82378 68886
rect 94826 68838 94862 77189
rect 94910 77169 94946 77174
rect 94902 77163 94954 77169
rect 94902 77105 94954 77111
rect 82426 68802 94862 68838
rect 82334 12462 82386 12468
rect 82334 12404 82386 12410
rect 82342 12400 82378 12404
rect 82426 12384 82462 68802
rect 94910 68754 94946 77105
rect 94994 77085 95030 77090
rect 94986 77079 95038 77085
rect 94986 77021 95038 77027
rect 82510 68718 94946 68754
rect 82418 12378 82470 12384
rect 82418 12320 82470 12326
rect 82426 12316 82462 12320
rect 82510 12300 82546 68718
rect 94994 68670 95030 77021
rect 95078 77001 95114 77006
rect 95070 76995 95122 77001
rect 95070 76937 95122 76943
rect 82594 68634 95030 68670
rect 82502 12294 82554 12300
rect 82502 12236 82554 12242
rect 82510 12232 82546 12236
rect 82594 12216 82630 68634
rect 95078 68586 95114 76937
rect 95162 76917 95198 76922
rect 95154 76911 95206 76917
rect 95154 76853 95206 76859
rect 82678 68550 95114 68586
rect 82586 12210 82638 12216
rect 82586 12152 82638 12158
rect 82594 12148 82630 12152
rect 82678 12132 82714 68550
rect 95162 68502 95198 76853
rect 95246 76833 95282 76838
rect 95238 76827 95290 76833
rect 95238 76769 95290 76775
rect 82762 68466 95198 68502
rect 82670 12126 82722 12132
rect 82670 12068 82722 12074
rect 82678 12064 82714 12068
rect 82762 12048 82798 68466
rect 95246 68418 95282 76769
rect 95330 76749 95366 76754
rect 95322 76743 95374 76749
rect 95322 76685 95374 76691
rect 82846 68382 95282 68418
rect 82754 12042 82806 12048
rect 82754 11984 82806 11990
rect 82762 11980 82798 11984
rect 82846 11964 82882 68382
rect 95330 68334 95366 76685
rect 95414 76665 95450 76670
rect 95406 76659 95458 76665
rect 95406 76601 95458 76607
rect 82930 68298 95366 68334
rect 82838 11958 82890 11964
rect 82838 11900 82890 11906
rect 82846 11896 82882 11900
rect 82930 11880 82966 68298
rect 95414 68250 95450 76601
rect 95498 76581 95534 76586
rect 95490 76575 95542 76581
rect 95490 76517 95542 76523
rect 83014 68214 95450 68250
rect 82922 11874 82974 11880
rect 82922 11816 82974 11822
rect 82930 11812 82966 11816
rect 83014 11796 83050 68214
rect 95498 68166 95534 76517
rect 143503 75327 143553 78351
rect 143502 75321 143554 75327
rect 143502 75263 143554 75269
rect 147356 71047 147520 80966
rect 147658 80966 148622 81390
rect 147658 75178 147822 80966
rect 151999 80962 153147 81394
rect 147921 75414 147971 78352
rect 151999 75690 152140 80962
rect 156819 79797 157122 81513
rect 152455 75586 152505 78348
rect 158308 77961 158344 89591
rect 160429 82089 160805 82143
rect 160429 80742 160460 82089
rect 160761 80742 160805 82089
rect 160429 80685 160805 80742
rect 160959 81841 161338 81881
rect 160959 80732 160996 81841
rect 161307 80732 161338 81841
rect 160959 80688 161338 80732
rect 176097 80169 176409 88365
rect 178193 80169 178505 88328
rect 193813 82259 194192 82310
rect 193282 81893 193664 81934
rect 193282 81115 193329 81893
rect 193632 81115 193664 81893
rect 193282 81070 193664 81115
rect 193813 81115 193852 82259
rect 194157 81115 194192 82259
rect 193813 81076 194192 81115
rect 196230 78044 196266 89828
rect 196538 83144 196716 96865
rect 262998 95385 263296 111182
rect 263932 98918 264232 113136
rect 264754 103448 265082 111968
rect 265604 106856 265914 113535
rect 267203 108437 267209 108489
rect 267261 108437 267267 108489
rect 267089 108417 267141 108423
rect 267089 108359 267141 108365
rect 267219 108359 267252 108437
rect 266973 108351 267005 108359
rect 266964 108345 267016 108351
rect 266964 108287 267016 108293
rect 266840 108273 266892 108280
rect 266973 108279 267006 108287
rect 266840 108215 266892 108221
rect 266850 107877 266882 108215
rect 266974 108202 267006 108279
rect 266840 107871 266892 107877
rect 266973 107874 267005 108202
rect 266840 107813 266892 107819
rect 266963 107868 267015 107874
rect 267095 107854 267127 108359
rect 267220 107870 267252 108359
rect 272872 108201 272924 108207
rect 272872 108143 272924 108149
rect 272747 108129 272799 108135
rect 272747 108071 272799 108077
rect 272757 107898 272789 108071
rect 272882 107907 272914 108143
rect 272872 107901 272924 107907
rect 272747 107892 272799 107898
rect 267210 107864 267262 107870
rect 266963 107810 267015 107816
rect 267079 107802 267085 107854
rect 267137 107802 267143 107854
rect 272872 107843 272924 107849
rect 272747 107834 272799 107840
rect 267210 107806 267262 107812
rect 265604 106546 266264 106856
rect 278768 106796 279036 114000
rect 278416 106528 279036 106796
rect 264754 103120 266350 103448
rect 279583 103348 279893 110110
rect 278458 103038 279893 103348
rect 263932 98618 266294 98918
rect 280295 98744 280585 114394
rect 278458 98454 280585 98744
rect 262998 95087 266313 95385
rect 281112 95274 281380 110728
rect 293208 108400 293454 111316
rect 293808 108400 294054 112604
rect 299130 108376 299376 110052
rect 299730 108376 299976 111960
rect 305052 108440 305298 109396
rect 305664 108440 305910 110698
rect 286469 103061 286531 103067
rect 286469 102993 286531 102999
rect 286389 102768 286441 102774
rect 286389 102710 286441 102716
rect 278478 95006 281380 95274
rect 198816 90609 200405 90631
rect 198816 90469 198858 90609
rect 200372 90469 200405 90609
rect 198816 90451 200405 90469
rect 198814 89070 200403 89092
rect 198814 88930 198845 89070
rect 200359 88930 200403 89070
rect 198814 88912 200403 88930
rect 196538 83143 207806 83144
rect 196538 82881 207863 83143
rect 196538 82880 196716 82881
rect 207615 82094 207863 82881
rect 198378 81660 199826 82084
rect 202733 81660 204237 82087
rect 207615 81662 208688 82094
rect 198378 79784 198678 81660
rect 202730 81098 203106 81530
rect 207241 81101 207566 81525
rect 163169 78038 163221 78044
rect 196222 78038 196274 78044
rect 191480 78030 191486 78038
rect 163221 77994 191486 78030
rect 191480 77986 191486 77994
rect 191538 77986 191544 78038
rect 163169 77980 163221 77986
rect 196222 77980 196274 77986
rect 158300 77955 158352 77961
rect 158300 77897 158352 77903
rect 158308 77894 158344 77897
rect 199065 76004 199115 78491
rect 199064 75998 199116 76004
rect 199064 75940 199116 75946
rect 152454 75580 152506 75586
rect 152454 75522 152506 75528
rect 147920 75408 147972 75414
rect 147920 75350 147972 75356
rect 202942 70536 203106 81098
rect 203483 75837 203533 78489
rect 203482 75831 203534 75837
rect 203482 75773 203534 75779
rect 207402 70023 207566 81101
rect 207730 81101 208697 81525
rect 207730 72071 207894 81101
rect 208017 75749 208067 78475
rect 208016 75743 208068 75749
rect 208016 75685 208068 75691
rect 83098 68130 95534 68166
rect 83006 11790 83058 11796
rect 83006 11732 83058 11738
rect 83014 11728 83050 11732
rect 83098 11712 83134 68130
rect 83665 61969 83739 61975
rect 83298 58821 83334 58832
rect 83288 58815 83340 58821
rect 83288 58757 83340 58763
rect 83090 11706 83142 11712
rect 83090 11648 83142 11654
rect 81705 10874 81757 10880
rect 81705 10816 81757 10822
rect 81713 10811 81749 10816
rect 35520 5854 35572 5860
rect 35520 5796 35572 5802
rect 35528 5792 35564 5796
rect 83298 2775 83334 58757
rect 83382 52554 83418 52558
rect 83370 52548 83422 52554
rect 83370 52490 83422 52496
rect 83290 2769 83342 2775
rect 83290 2711 83342 2717
rect 83298 2706 83334 2711
rect 83382 2691 83418 52490
rect 83466 46903 83502 46910
rect 83460 46897 83512 46903
rect 83460 46839 83512 46845
rect 83374 2685 83426 2691
rect 83374 2627 83426 2633
rect 83382 2624 83418 2627
rect 83466 2607 83502 46839
rect 83550 40636 83586 40642
rect 83546 40630 83598 40636
rect 83546 40572 83598 40578
rect 83458 2601 83510 2607
rect 83458 2543 83510 2549
rect 83466 2538 83502 2543
rect 83550 2523 83586 40572
rect 83665 2611 83739 61744
rect 83832 28201 84087 65026
rect 84254 61958 84306 61964
rect 84254 61900 84306 61906
rect 84262 60430 84298 61900
rect 84262 60394 86046 60430
rect 84262 48520 84298 60394
rect 84763 59287 86016 59309
rect 84763 58525 84783 59287
rect 84916 59257 86016 59287
rect 84916 59072 84944 59257
rect 84916 59020 86016 59072
rect 84916 58561 84944 59020
rect 84916 58525 86016 58561
rect 84763 58509 86016 58525
rect 84766 51474 86016 51492
rect 84766 50906 84782 51474
rect 84925 51440 86016 51474
rect 84925 51152 84941 51440
rect 84925 51100 86016 51152
rect 84925 50940 84941 51100
rect 84925 50906 86016 50940
rect 84766 50888 86016 50906
rect 84766 50887 84941 50888
rect 84262 48484 86030 48520
rect 84829 47391 84838 47395
rect 84802 47339 84838 47391
rect 84829 47335 84838 47339
rect 84898 47391 84907 47395
rect 84898 47339 86018 47391
rect 84898 47335 84907 47339
rect 84827 47154 84836 47158
rect 84802 47102 84836 47154
rect 84827 47098 84836 47102
rect 84896 47154 84905 47158
rect 84896 47102 86018 47154
rect 84896 47098 84905 47102
rect 84827 46643 84836 46647
rect 84808 46591 84836 46643
rect 84827 46587 84836 46591
rect 84896 46643 84905 46647
rect 84896 46591 86020 46643
rect 84896 46587 84905 46591
rect 84797 39574 84806 39578
rect 84786 39522 84806 39574
rect 84797 39518 84806 39522
rect 84866 39574 84875 39578
rect 84866 39522 86020 39574
rect 84866 39518 84875 39522
rect 84801 39234 84810 39238
rect 84786 39182 84810 39234
rect 84801 39178 84810 39182
rect 84870 39234 84879 39238
rect 84870 39182 86020 39234
rect 84870 39178 84879 39182
rect 84797 39022 84806 39026
rect 84786 38970 84806 39022
rect 84797 38966 84806 38970
rect 84866 39022 84875 39026
rect 84866 38970 86020 39022
rect 84866 38966 84875 38970
rect 131043 28201 131298 65539
rect 133981 34870 134181 66026
rect 134730 60170 134938 69605
rect 134361 59962 134938 60170
rect 134361 48217 134569 59962
rect 170105 58888 170252 63473
rect 183932 59797 185250 59846
rect 183932 59273 183998 59797
rect 185192 59273 185250 59797
rect 183932 59224 185250 59273
rect 186053 54394 186170 61704
rect 189741 58513 190803 58535
rect 186821 57945 186969 58457
rect 189741 58319 189798 58513
rect 190768 58319 190803 58513
rect 189741 58275 190803 58319
rect 186821 57797 187456 57945
rect 191384 56017 191523 64524
rect 190840 55878 191523 56017
rect 186822 55305 187400 55431
rect 186242 54020 186294 54027
rect 186242 53962 186294 53968
rect 182377 52696 184035 52741
rect 182377 52513 182438 52696
rect 183994 52513 184035 52696
rect 182377 52464 184035 52513
rect 186250 48685 186286 53962
rect 186822 53484 186948 55305
rect 191072 55017 192134 55048
rect 191072 55012 191120 55017
rect 190678 54832 191120 55012
rect 192099 54832 192134 55017
rect 190678 54818 192134 54832
rect 191072 54788 192134 54818
rect 186469 52604 187820 52655
rect 186469 52451 186566 52604
rect 186479 52384 186566 52451
rect 187774 52384 187820 52604
rect 186479 52333 187820 52384
rect 186250 48649 189261 48685
rect 134361 47905 134394 48217
rect 134530 47905 134569 48217
rect 134361 47893 134569 47905
rect 133981 34558 134004 34870
rect 134140 34558 134181 34870
rect 133981 34549 134181 34558
rect 186255 34827 188561 34858
rect 186255 34181 186599 34827
rect 188523 34181 188561 34827
rect 186255 34150 188561 34181
rect 174601 33529 175385 33629
rect 174601 33169 175434 33269
rect 175028 31631 176381 31682
rect 175028 31064 175103 31631
rect 176317 31064 176381 31631
rect 175028 30976 176381 31064
rect 83832 27946 84384 28201
rect 130679 27946 131298 28201
rect 174703 30337 175796 30437
rect 173960 27930 173996 27950
rect 173952 27924 174004 27930
rect 173952 27866 174004 27872
rect 124105 12624 124487 12672
rect 90535 12520 90924 12560
rect 90535 10985 90573 12520
rect 90888 10985 90924 12520
rect 123574 11829 123957 11867
rect 90535 10924 90924 10985
rect 91072 11779 91458 11822
rect 91072 10993 91116 11779
rect 91423 10993 91458 11779
rect 91072 10933 91458 10993
rect 92028 10982 92080 10988
rect 92028 10924 92080 10930
rect 93466 10982 93518 10988
rect 93466 10924 93518 10930
rect 95094 10982 95146 10988
rect 95094 10924 95146 10930
rect 96722 10982 96774 10988
rect 96722 10924 96774 10930
rect 98350 10982 98402 10988
rect 98350 10924 98402 10930
rect 99978 10982 100030 10988
rect 99978 10924 100030 10930
rect 101606 10982 101658 10988
rect 101606 10924 101658 10930
rect 103234 10982 103286 10988
rect 103234 10924 103286 10930
rect 104862 10982 104914 10988
rect 104862 10924 104914 10930
rect 110099 10986 110174 10996
rect 110099 10928 110109 10986
rect 110167 10928 110174 10986
rect 92036 9704 92072 10924
rect 92028 9698 92080 9704
rect 92028 9640 92080 9646
rect 93474 9284 93510 10924
rect 93466 9278 93518 9284
rect 93466 9220 93518 9226
rect 95102 9201 95138 10924
rect 95094 9195 95146 9201
rect 95094 9137 95146 9143
rect 96730 9113 96766 10924
rect 96722 9107 96774 9113
rect 96722 9049 96774 9055
rect 98358 9029 98394 10924
rect 98350 9023 98402 9029
rect 98350 8965 98402 8971
rect 99986 8945 100022 10924
rect 99978 8939 100030 8945
rect 99978 8881 100030 8887
rect 101614 8861 101650 10924
rect 101606 8855 101658 8861
rect 101606 8797 101658 8803
rect 103242 8777 103278 10924
rect 103234 8771 103286 8777
rect 103234 8713 103286 8719
rect 104870 8699 104906 10924
rect 110099 10921 110174 10928
rect 111727 10986 111802 10996
rect 111727 10928 111737 10986
rect 111795 10928 111802 10986
rect 111727 10921 111802 10928
rect 113355 10986 113430 10996
rect 113355 10928 113365 10986
rect 113423 10928 113430 10986
rect 113355 10921 113430 10928
rect 114983 10986 115058 10996
rect 114983 10928 114993 10986
rect 115051 10928 115058 10986
rect 114983 10921 115058 10928
rect 116611 10986 116686 10996
rect 116611 10928 116621 10986
rect 116679 10928 116686 10986
rect 116611 10921 116686 10928
rect 118239 10986 118314 10996
rect 118239 10928 118249 10986
rect 118307 10928 118314 10986
rect 118239 10921 118314 10928
rect 119867 10986 119942 10996
rect 119867 10928 119877 10986
rect 119935 10928 119942 10986
rect 119867 10921 119942 10928
rect 121494 10986 121569 10995
rect 121494 10928 121505 10986
rect 121563 10928 121569 10986
rect 123574 10977 123624 11829
rect 123927 10977 123957 11829
rect 123574 10929 123957 10977
rect 124105 10975 124147 12624
rect 124449 10975 124487 12624
rect 124105 10928 124487 10975
rect 110112 9791 110155 10921
rect 111740 9876 111783 10921
rect 113368 9956 113411 10921
rect 114996 10046 115039 10921
rect 116624 10125 116667 10921
rect 118252 10213 118295 10921
rect 119877 10287 119935 10921
rect 121494 10920 121569 10928
rect 121505 10377 121563 10920
rect 121505 10313 121563 10319
rect 119877 10223 119935 10229
rect 118248 10207 118300 10213
rect 118248 10149 118300 10155
rect 116620 10119 116672 10125
rect 116620 10061 116672 10067
rect 114992 10040 115044 10046
rect 114992 9982 115044 9988
rect 113358 9904 113364 9956
rect 113416 9904 113422 9956
rect 111736 9870 111788 9876
rect 111736 9812 111788 9818
rect 110108 9785 110160 9791
rect 110108 9727 110160 9733
rect 104862 8693 104914 8699
rect 104862 8635 104914 8641
rect 173960 8528 173996 27866
rect 83542 2517 83594 2523
rect 83542 2459 83594 2465
rect 83550 2449 83586 2459
rect 31561 2411 31835 2418
rect 31561 2330 31835 2337
rect 83665 2331 83739 2337
rect 31561 0 31631 2330
rect 135662 1935 135698 7929
rect 135654 1929 135706 1935
rect 135654 1871 135706 1877
rect 138118 1850 138154 7961
rect 140624 6269 140652 7925
rect 143133 6449 143161 7940
rect 145606 6599 145634 7937
rect 148195 6725 148223 7937
rect 150580 6880 150608 7955
rect 153150 7671 153178 7948
rect 152368 7643 153178 7671
rect 150580 6852 152284 6880
rect 148195 6697 152172 6725
rect 145606 6571 152060 6599
rect 143133 6421 151948 6449
rect 140624 6241 151836 6269
rect 138110 1844 138162 1850
rect 138110 1786 138162 1792
rect 151808 0 151836 6241
rect 151920 0 151948 6421
rect 152032 0 152060 6571
rect 152144 0 152172 6697
rect 152256 0 152284 6852
rect 152368 0 152396 7643
rect 155630 7512 155658 7957
rect 152480 7484 155658 7512
rect 152480 0 152508 7484
rect 158114 7331 158142 7935
rect 152592 7303 158142 7331
rect 152592 0 152620 7303
rect 152704 7193 152732 7198
rect 160622 7193 160650 7980
rect 152704 7165 160650 7193
rect 152704 0 152732 7165
rect 163125 7013 163153 7957
rect 152816 6985 163153 7013
rect 152816 0 152844 6985
rect 165631 6870 165659 7965
rect 152928 6842 165659 6870
rect 152928 0 152956 6842
rect 168117 6684 168145 7944
rect 173952 7782 174004 8528
rect 173952 7723 174004 7730
rect 153040 6656 168145 6684
rect 153040 0 153068 6656
rect 153152 0 153180 6269
rect 153264 0 153292 6269
rect 153376 0 153404 6269
rect 153488 0 153516 6269
rect 174703 1996 174803 30337
rect 175029 29713 176382 29766
rect 175029 29146 175090 29713
rect 176304 29146 176382 29713
rect 175029 29060 176382 29146
rect 186616 28994 188515 28995
rect 186283 28962 188515 28994
rect 186283 28312 186663 28962
rect 188472 28312 188515 28962
rect 186283 28286 188515 28312
rect 186616 28284 188515 28286
rect 174703 1804 174729 1996
rect 174781 1804 174803 1996
rect 174703 1794 174803 1804
rect 189225 1767 189261 48649
rect 192668 34679 192868 66563
rect 193326 48053 193499 69006
rect 214920 66004 215276 78748
rect 215384 75158 215420 78457
rect 215376 75152 215428 75158
rect 215376 75094 215428 75100
rect 219436 72150 219792 78748
rect 219900 75918 219936 78455
rect 219892 75912 219944 75918
rect 219892 75854 219944 75860
rect 223952 71134 224308 78806
rect 224416 75496 224452 78444
rect 224408 75490 224460 75496
rect 224408 75432 224460 75438
rect 228657 64906 229087 78470
rect 230711 65446 231141 78454
rect 231386 76082 231422 78446
rect 231378 76076 231430 76082
rect 231378 76018 231430 76024
rect 235384 72596 235740 78778
rect 235902 75666 235938 78475
rect 235894 75660 235946 75666
rect 235894 75602 235946 75608
rect 239900 71536 240256 78746
rect 240418 75241 240454 78448
rect 240410 75235 240462 75241
rect 240410 75177 240462 75183
rect 229065 58888 229212 63999
rect 237206 60562 237342 65580
rect 241322 60594 241458 65074
rect 241722 60594 241858 66612
rect 244416 66446 244772 78746
rect 281972 75840 282108 75848
rect 277831 75150 277986 75200
rect 245838 60660 245974 66102
rect 246238 60660 246374 67542
rect 250354 60628 250490 67135
rect 250754 60628 250890 68638
rect 254870 60628 255006 68149
rect 255270 60628 255406 70188
rect 259386 60660 259522 70718
rect 259786 60660 259922 72250
rect 263902 60660 264038 72754
rect 264302 60660 264438 71228
rect 268418 60660 268554 71736
rect 268818 60660 268954 74300
rect 272934 60628 273070 74796
rect 273334 60628 273470 73280
rect 277450 60660 277586 73794
rect 277850 60660 277986 75150
rect 281972 60572 282108 75712
rect 241188 51074 241216 52179
rect 249601 52167 249653 52173
rect 241522 51363 241550 52147
rect 241606 51633 241634 52134
rect 241594 51627 241646 51633
rect 241594 51569 241646 51575
rect 241907 51490 241935 52158
rect 241895 51484 241947 51490
rect 241895 51426 241947 51432
rect 241510 51357 241562 51363
rect 241510 51299 241562 51305
rect 246027 51198 246063 52157
rect 249601 52109 249653 52115
rect 248173 52008 248225 52014
rect 248173 51950 248225 51956
rect 246019 51192 246071 51198
rect 246019 51134 246071 51140
rect 248007 51192 248059 51198
rect 248007 51134 248059 51140
rect 241170 51022 241176 51074
rect 241228 51022 241234 51074
rect 243689 34975 246588 35026
rect 243689 34357 244169 34975
rect 246537 34357 246588 34975
rect 243689 34318 246588 34357
rect 231789 33676 232852 33776
rect 231789 33316 232854 33416
rect 232626 31763 234573 31847
rect 232626 31208 232705 31763
rect 234494 31208 234573 31763
rect 232626 31141 234573 31208
rect 232269 30511 233250 30611
rect 232269 29934 232369 30511
rect 232269 29228 232370 29934
rect 232627 29867 234573 29934
rect 232627 29312 232969 29867
rect 234511 29312 234573 29867
rect 232627 29228 234573 29312
rect 194601 2187 194637 8101
rect 194593 2181 194645 2187
rect 194593 2123 194645 2129
rect 197084 2102 197120 8067
rect 199592 6168 199620 8099
rect 202092 6267 202120 8085
rect 204548 6445 204576 8074
rect 207041 6582 207069 8089
rect 209599 7818 209627 8109
rect 209599 7790 211076 7818
rect 207041 6554 210964 6582
rect 204548 6417 210852 6445
rect 202092 6239 210740 6267
rect 210600 6168 210628 6169
rect 199592 6140 210628 6168
rect 197076 2096 197128 2102
rect 197076 2038 197128 2044
rect 189217 1761 189269 1767
rect 189217 1703 189269 1709
rect 210600 0 210628 6140
rect 210712 0 210740 6239
rect 210824 0 210852 6417
rect 210936 0 210964 6554
rect 211048 0 211076 7790
rect 212110 7672 212138 8076
rect 211160 7644 212138 7672
rect 211160 0 211188 7644
rect 214572 7474 214600 8107
rect 211272 7446 214600 7474
rect 211272 0 211300 7446
rect 217069 7324 217097 8093
rect 211384 7296 217097 7324
rect 211384 0 211412 7296
rect 219585 7149 219613 8080
rect 211496 7121 219613 7149
rect 211496 0 211524 7121
rect 222077 6951 222105 8103
rect 211608 6923 222105 6951
rect 211608 0 211636 6923
rect 224567 6756 224595 8120
rect 211720 6728 224595 6756
rect 211720 0 211748 6728
rect 227053 6595 227081 8062
rect 211832 6567 227081 6595
rect 211832 0 211860 6567
rect 211944 0 211972 6169
rect 212056 0 212084 6169
rect 212168 0 212196 6169
rect 212280 0 212308 6169
rect 232269 2265 232369 29228
rect 243716 29128 247186 29162
rect 243716 28490 244399 29128
rect 247152 28490 247186 29128
rect 243716 28454 247186 28490
rect 233042 28384 233094 28390
rect 233042 28326 233094 28332
rect 233050 7872 233086 28326
rect 233042 7866 233094 7872
rect 233042 7808 233094 7814
rect 248013 4732 248049 51134
rect 248097 47551 248133 47561
rect 248082 47545 248134 47551
rect 248082 47487 248134 47493
rect 248005 4726 248057 4732
rect 248005 4668 248057 4674
rect 248097 4648 248133 47487
rect 248089 4642 248141 4648
rect 248089 4584 248141 4590
rect 248181 4564 248217 51950
rect 248677 51918 248729 51924
rect 248677 51860 248729 51866
rect 248265 42918 248301 42920
rect 248259 42912 248311 42918
rect 248259 42854 248311 42860
rect 248173 4558 248225 4564
rect 248173 4500 248225 4506
rect 248265 4480 248301 42854
rect 248257 4474 248309 4480
rect 248257 4416 248309 4422
rect 248685 4060 248721 51860
rect 249433 51838 249485 51844
rect 249433 51780 249485 51786
rect 248937 51719 248973 51736
rect 248929 51713 248981 51719
rect 248929 51655 248981 51661
rect 248769 42834 248805 42836
rect 248758 42828 248810 42834
rect 248758 42770 248810 42776
rect 248677 4054 248729 4060
rect 248677 3996 248729 4002
rect 248769 3976 248805 42770
rect 248761 3970 248813 3976
rect 248761 3912 248813 3918
rect 248937 3808 248973 51655
rect 249009 47461 249061 47467
rect 249009 47403 249061 47409
rect 248929 3802 248981 3808
rect 248929 3744 248981 3750
rect 249021 3724 249057 47403
rect 249013 3718 249065 3724
rect 249013 3660 249065 3666
rect 249441 3304 249477 51780
rect 249515 42744 249567 42750
rect 249515 42686 249567 42692
rect 249433 3298 249485 3304
rect 249433 3240 249485 3246
rect 249525 3220 249561 42686
rect 249517 3214 249569 3220
rect 249517 3156 249569 3162
rect 249609 3136 249645 52109
rect 250555 51723 250591 52140
rect 250547 51717 250599 51723
rect 250547 51659 250599 51665
rect 249769 51627 249821 51633
rect 249769 51569 249821 51575
rect 249687 47377 249739 47383
rect 249687 47319 249739 47325
rect 249601 3130 249653 3136
rect 249601 3072 249653 3078
rect 249693 3052 249729 47319
rect 249685 3046 249737 3052
rect 249685 2988 249737 2994
rect 249777 2969 249813 51569
rect 249853 51488 249905 51494
rect 249853 51430 249905 51436
rect 249769 2963 249821 2969
rect 249769 2905 249821 2911
rect 249861 2885 249897 51430
rect 249937 51354 249989 51360
rect 249937 51296 249989 51302
rect 249853 2879 249905 2885
rect 249853 2821 249905 2827
rect 249945 2800 249981 51296
rect 250029 51080 250065 51090
rect 250022 51074 250074 51080
rect 250022 51016 250074 51022
rect 249937 2794 249989 2800
rect 249937 2736 249989 2742
rect 250029 2716 250065 51016
rect 276858 32206 277828 32722
rect 280310 32222 281280 32738
rect 273484 31314 273536 31320
rect 273484 31256 273536 31262
rect 273408 31199 273444 31208
rect 273400 31193 273452 31199
rect 273400 31135 273452 31141
rect 257238 26004 257390 26022
rect 257238 24982 257258 26004
rect 257372 24982 257390 26004
rect 257238 24958 257390 24982
rect 250021 2710 250073 2716
rect 250021 2652 250073 2658
rect 232269 2073 232290 2265
rect 232342 2073 232369 2265
rect 232269 2055 232369 2073
rect 255683 463 255775 24008
rect 256055 790 256147 23821
rect 273408 1684 273444 31135
rect 273400 1678 273452 1684
rect 273400 1620 273452 1626
rect 273408 1617 273444 1620
rect 273492 1600 273528 31256
rect 273660 25413 273696 25425
rect 273652 25407 273704 25413
rect 273652 25349 273704 25355
rect 273576 25292 273612 25307
rect 273568 25286 273620 25292
rect 273568 25228 273620 25234
rect 273484 1594 273536 1600
rect 273484 1536 273536 1542
rect 273492 1532 273528 1536
rect 273576 1516 273612 25228
rect 273568 1510 273620 1516
rect 273568 1452 273620 1458
rect 273576 1447 273612 1452
rect 273660 1432 273696 25349
rect 276858 19302 277830 19838
rect 280310 19302 281282 19838
rect 286397 2632 286433 102710
rect 286389 2626 286441 2632
rect 286389 2568 286441 2574
rect 286481 2549 286517 102993
rect 287314 101176 287366 101182
rect 287314 101118 287366 101124
rect 287230 101092 287282 101098
rect 287230 101034 287282 101040
rect 287061 100841 287113 100847
rect 287061 100783 287113 100789
rect 286893 93305 286945 93311
rect 286893 93247 286945 93253
rect 286649 87012 286685 87014
rect 286636 87006 286696 87012
rect 286636 86940 286696 86946
rect 286557 86702 286609 86708
rect 286557 86644 286609 86650
rect 286473 2543 286525 2549
rect 286473 2485 286525 2491
rect 286565 2464 286601 86644
rect 286557 2458 286609 2464
rect 286557 2400 286609 2406
rect 286649 2381 286685 86940
rect 286810 85100 286862 85106
rect 286810 85042 286862 85048
rect 286725 85016 286777 85022
rect 286725 84958 286777 84964
rect 286733 5068 286769 84958
rect 286725 5062 286777 5068
rect 286725 5004 286777 5010
rect 286817 4984 286853 85042
rect 286901 82756 286937 93247
rect 286985 93230 287021 93231
rect 286977 93224 287029 93230
rect 286977 93166 287029 93172
rect 286985 82840 287021 93166
rect 287069 85423 287105 100783
rect 287153 100762 287189 100764
rect 287145 100756 287197 100762
rect 287145 100698 287197 100704
rect 287153 85500 287189 100698
rect 287237 85578 287273 101034
rect 287321 85659 287357 101118
rect 287741 101015 287777 101023
rect 287733 101009 287785 101015
rect 287733 100951 287785 100957
rect 287480 93138 287532 93144
rect 287480 93080 287532 93086
rect 287398 93054 287450 93060
rect 287398 92996 287450 93002
rect 287405 85751 287441 92996
rect 287489 85831 287525 93080
rect 287565 92969 287617 92975
rect 287565 92911 287617 92917
rect 287573 85913 287609 92911
rect 287649 92888 287701 92894
rect 287649 92830 287701 92836
rect 287657 85986 287693 92830
rect 287741 86086 287777 100951
rect 287825 100933 287861 100937
rect 287817 100927 287869 100933
rect 287817 100869 287869 100875
rect 287825 86188 287861 100869
rect 311675 95024 311905 111346
rect 312366 98524 312566 114730
rect 313038 103228 313288 111970
rect 314180 106624 314380 114240
rect 321596 109428 321648 109434
rect 321596 109370 321648 109376
rect 321350 109188 321402 109194
rect 321350 109130 321402 109136
rect 315446 108948 315498 108954
rect 315446 108890 315498 108896
rect 315452 107768 315492 108890
rect 315558 108828 315610 108834
rect 315558 108770 315610 108776
rect 315562 107778 315602 108770
rect 315678 108708 315730 108714
rect 315678 108650 315730 108656
rect 315684 107792 315724 108650
rect 315804 108588 315856 108594
rect 315804 108530 315856 108536
rect 315810 107792 315850 108530
rect 321356 107944 321396 109130
rect 321468 109068 321520 109074
rect 321468 109010 321520 109016
rect 321474 107944 321514 109010
rect 321602 107954 321642 109370
rect 321718 109308 321770 109314
rect 321718 109250 321770 109256
rect 321596 107948 321648 107954
rect 321724 107950 321764 109250
rect 321350 107938 321402 107944
rect 321350 107880 321402 107886
rect 321468 107938 321520 107944
rect 321712 107898 321718 107950
rect 321770 107898 321776 107950
rect 321596 107890 321648 107896
rect 321468 107880 321520 107886
rect 315678 107786 315730 107792
rect 315556 107772 315608 107778
rect 315446 107762 315498 107768
rect 315678 107728 315730 107734
rect 315804 107786 315856 107792
rect 315804 107728 315856 107734
rect 315556 107714 315608 107720
rect 315446 107704 315498 107710
rect 314180 106424 314878 106624
rect 327454 106594 327654 113646
rect 327006 106394 327654 106594
rect 313038 102978 314978 103228
rect 328007 103062 328237 110128
rect 327054 102832 328237 103062
rect 329106 98610 329306 113210
rect 312366 98324 314868 98524
rect 326954 98410 329306 98610
rect 329830 95108 330102 110754
rect 360457 107582 361047 111805
rect 410154 105365 410444 111889
rect 412615 105311 412903 111358
rect 463511 107592 464085 111274
rect 412749 105303 412903 105311
rect 311675 94794 314914 95024
rect 327096 94836 330102 95108
rect 388877 90856 390307 90889
rect 388877 90725 388908 90856
rect 390258 90725 390307 90856
rect 388877 90694 390307 90725
rect 388959 89308 390389 89349
rect 388959 89177 388995 89308
rect 390345 89177 390389 89308
rect 388959 89154 390389 89177
rect 287825 86152 288029 86188
rect 287741 86050 287945 86086
rect 287657 85950 287861 85986
rect 287573 85877 287777 85913
rect 287489 85795 287693 85831
rect 287405 85715 287609 85751
rect 287321 85658 287520 85659
rect 287321 85623 287525 85658
rect 287237 85542 287441 85578
rect 287153 85464 287357 85500
rect 287069 85387 287273 85423
rect 287146 84932 287198 84938
rect 287146 84874 287198 84880
rect 287062 84848 287114 84854
rect 287062 84790 287114 84796
rect 286977 82834 287029 82840
rect 286977 82776 287029 82782
rect 286893 82750 286945 82756
rect 286893 82692 286945 82698
rect 286978 77062 287030 77068
rect 286978 77004 287030 77010
rect 286894 76978 286946 76984
rect 286894 76920 286946 76926
rect 286809 4978 286861 4984
rect 286809 4920 286861 4926
rect 286901 4900 286937 76920
rect 286893 4894 286945 4900
rect 286893 4836 286945 4842
rect 286985 4816 287021 77004
rect 286977 4810 287029 4816
rect 286977 4752 287029 4758
rect 287069 4396 287105 84790
rect 287061 4390 287113 4396
rect 287061 4332 287113 4338
rect 287153 4312 287189 84874
rect 287237 82923 287273 85387
rect 287321 83007 287357 85464
rect 287313 83001 287365 83007
rect 287313 82943 287365 82949
rect 287229 82917 287281 82923
rect 287229 82859 287281 82865
rect 287312 76894 287364 76900
rect 287312 76836 287364 76842
rect 287229 76810 287281 76816
rect 287229 76752 287281 76758
rect 287145 4306 287197 4312
rect 287145 4248 287197 4254
rect 287237 4228 287273 76752
rect 287229 4222 287281 4228
rect 287229 4164 287281 4170
rect 287321 4144 287357 76836
rect 287313 4138 287365 4144
rect 287313 4080 287365 4086
rect 287405 3640 287441 85542
rect 287397 3634 287449 3640
rect 287397 3576 287449 3582
rect 287489 3556 287525 85623
rect 287481 3550 287533 3556
rect 287481 3492 287533 3498
rect 287573 3472 287609 85715
rect 287565 3466 287617 3472
rect 287565 3408 287617 3414
rect 287657 3388 287693 85795
rect 287741 83090 287777 85877
rect 287825 83174 287861 85950
rect 287909 83258 287945 86050
rect 287993 83342 288029 86152
rect 289605 84764 289657 84770
rect 289605 84706 289657 84712
rect 287985 83336 288037 83342
rect 287985 83278 288037 83284
rect 289017 83338 289069 83344
rect 289017 83280 289069 83286
rect 287901 83252 287953 83258
rect 287901 83194 287953 83200
rect 288933 83254 288985 83260
rect 288933 83196 288985 83202
rect 287817 83168 287869 83174
rect 287817 83110 287869 83116
rect 288849 83170 288901 83176
rect 288849 83112 288901 83118
rect 287733 83084 287785 83090
rect 287733 83026 287785 83032
rect 288765 83086 288817 83092
rect 288765 83028 288817 83034
rect 288345 83000 288397 83006
rect 288345 82942 288397 82948
rect 288261 82916 288313 82922
rect 288261 82858 288313 82864
rect 288185 82838 288221 82839
rect 288177 82832 288229 82838
rect 288177 82774 288229 82780
rect 288093 82748 288145 82754
rect 288093 82690 288145 82696
rect 288017 56817 288053 56843
rect 288010 56811 288062 56817
rect 288010 56753 288062 56759
rect 287849 52184 287885 52200
rect 287836 52178 287888 52184
rect 287836 52120 287888 52126
rect 287765 42918 287801 42936
rect 287764 42912 287816 42918
rect 287764 42854 287816 42860
rect 287649 3382 287701 3388
rect 287649 3324 287701 3330
rect 287765 3070 287801 42854
rect 287849 3154 287885 52120
rect 287933 47551 287969 47573
rect 287929 47545 287981 47551
rect 287929 47487 287981 47493
rect 287933 3238 287969 47487
rect 288017 3322 288053 56753
rect 288101 3406 288137 82690
rect 288185 3490 288221 82774
rect 288269 3574 288305 82858
rect 288353 3658 288389 82942
rect 288521 56733 288557 56744
rect 288510 56727 288562 56733
rect 288510 56669 288562 56675
rect 288437 47467 288473 47481
rect 288428 47461 288480 47467
rect 288428 47403 288480 47409
rect 288437 3742 288473 47403
rect 288521 3826 288557 56669
rect 288689 52100 288725 52108
rect 288684 52094 288736 52100
rect 288684 52036 288736 52042
rect 288605 42834 288641 42839
rect 288594 42828 288646 42834
rect 288594 42770 288646 42776
rect 288605 3910 288641 42770
rect 288689 3994 288725 52036
rect 288773 4078 288809 83028
rect 288857 4162 288893 83112
rect 288941 4246 288977 83196
rect 289025 4330 289061 83280
rect 289437 77230 289489 77236
rect 289437 77172 289489 77178
rect 289193 56649 289229 56666
rect 289188 56643 289240 56649
rect 289188 56585 289240 56591
rect 289109 47383 289145 47399
rect 289103 47377 289155 47383
rect 289103 47319 289155 47325
rect 289109 4414 289145 47319
rect 289193 4498 289229 56585
rect 289361 52016 289397 52034
rect 289356 52010 289408 52016
rect 289356 51952 289408 51958
rect 289277 42750 289313 42761
rect 289271 42744 289323 42750
rect 289271 42686 289323 42692
rect 289277 4582 289313 42686
rect 289361 4666 289397 51952
rect 289445 4750 289481 77172
rect 289529 77152 289565 77155
rect 289521 77146 289573 77152
rect 289521 77088 289573 77094
rect 289529 4834 289565 77088
rect 289613 4918 289649 84706
rect 289697 84685 289733 84687
rect 289689 84679 289741 84685
rect 289689 84621 289741 84627
rect 289697 5002 289733 84621
rect 392562 83383 392740 95599
rect 380263 83160 392740 83383
rect 380263 82081 380502 83160
rect 392562 83159 392740 83160
rect 394813 82606 395187 82661
rect 379903 81659 380502 82081
rect 379903 81657 380439 81659
rect 384421 81655 385955 82087
rect 388921 81648 389720 82075
rect 375653 81092 376853 81524
rect 379894 81098 379998 81520
rect 380338 81098 381376 81520
rect 370496 78188 370832 78193
rect 375653 74594 375817 81092
rect 380338 78566 380502 81098
rect 376249 78382 376299 78541
rect 378764 78402 380502 78566
rect 384847 81093 385879 81525
rect 376248 78376 376300 78382
rect 376248 78318 376300 78324
rect 378764 75280 378928 78402
rect 380667 78285 380717 78509
rect 380666 78279 380718 78285
rect 380666 78221 380718 78227
rect 384374 78188 384710 78193
rect 384847 75656 385011 81093
rect 389433 79413 389720 81648
rect 394813 80687 394851 82606
rect 395147 80687 395187 82606
rect 394813 80638 395187 80687
rect 395338 81462 395710 81521
rect 395338 80671 395370 81462
rect 395671 80671 395710 81462
rect 395338 80627 395710 80671
rect 410297 79769 410609 87965
rect 412393 79769 412705 87965
rect 430738 83354 430916 95539
rect 490571 95070 490805 111308
rect 491192 98536 491392 114524
rect 505217 113979 506392 114179
rect 492728 113398 492924 113756
rect 491813 103110 492047 111974
rect 492724 106610 492924 113398
rect 504656 110388 504708 110394
rect 504656 110330 504708 110336
rect 504536 110268 504588 110274
rect 504536 110210 504588 110216
rect 498988 109908 499040 109914
rect 498988 109850 499040 109856
rect 498876 109788 498928 109794
rect 498876 109730 498928 109736
rect 498746 109668 498798 109674
rect 498746 109610 498798 109616
rect 498626 109548 498678 109554
rect 498626 109490 498678 109496
rect 498632 107876 498672 109490
rect 498626 107870 498678 107876
rect 498752 107864 498792 109610
rect 498882 107866 498922 109730
rect 498626 107812 498678 107818
rect 498746 107858 498798 107864
rect 498746 107800 498798 107806
rect 498876 107860 498928 107866
rect 498994 107864 499034 109850
rect 498876 107802 498928 107808
rect 498988 107858 499040 107864
rect 504542 107860 504582 110210
rect 504662 107876 504702 110330
rect 504896 110148 504948 110154
rect 504896 110090 504948 110096
rect 504774 110028 504826 110034
rect 504774 109970 504826 109976
rect 504780 107888 504820 109970
rect 504774 107882 504826 107888
rect 504902 107886 504942 110090
rect 505217 108458 505417 113979
rect 505217 108258 506046 108458
rect 504656 107870 504708 107876
rect 504530 107808 504536 107860
rect 504588 107808 504594 107860
rect 504774 107824 504826 107830
rect 504896 107880 504948 107886
rect 504896 107822 504948 107828
rect 504656 107812 504708 107818
rect 498988 107800 499040 107806
rect 492724 106410 493280 106610
rect 505846 106532 506046 108258
rect 505512 106332 506046 106532
rect 491813 102876 493332 103110
rect 506278 102976 506478 110106
rect 505524 102776 506478 102976
rect 506771 98722 506971 113505
rect 507369 101649 507569 112578
rect 509019 107274 509025 107354
rect 509105 107334 509114 107354
rect 509105 107278 510793 107334
rect 509105 107274 509114 107278
rect 508920 104866 508926 104946
rect 509006 104938 509014 104946
rect 509006 104882 510759 104938
rect 509006 104866 509014 104882
rect 508824 102468 508830 102548
rect 508910 102542 508921 102548
rect 508910 102486 510764 102542
rect 508910 102468 508921 102486
rect 491192 98336 493420 98536
rect 506771 98504 506937 98722
rect 505420 98304 506937 98504
rect 490571 94836 493360 95070
rect 507368 94974 507568 101649
rect 508734 100088 508740 100168
rect 508820 100146 508829 100168
rect 508820 100090 510810 100146
rect 508820 100088 508829 100090
rect 508636 97672 508642 97752
rect 508722 97750 508733 97752
rect 508722 97694 510776 97750
rect 508722 97672 508733 97694
rect 551427 95957 551627 112955
rect 571528 112364 571568 112376
rect 571408 112244 571448 112270
rect 571288 112124 571328 112144
rect 571168 112004 571208 112024
rect 571048 111884 571088 111904
rect 570928 111764 570968 111770
rect 570808 111644 570848 111658
rect 570688 111524 570728 111546
rect 570568 111404 570608 111420
rect 570448 111284 570488 111314
rect 570328 111164 570368 111184
rect 570208 111044 570248 111064
rect 570088 110924 570128 110946
rect 569968 110804 570008 110826
rect 569848 110700 569888 110714
rect 569728 110574 569768 110580
rect 550875 95700 551627 95957
rect 509479 95282 509485 95362
rect 509565 95354 509576 95362
rect 509565 95298 510747 95354
rect 551840 95317 564013 95445
rect 509565 95282 509576 95298
rect 505540 94774 507568 94974
rect 509392 92892 509398 92972
rect 509478 92958 509487 92972
rect 509478 92902 510785 92958
rect 509478 92892 509487 92902
rect 434140 90895 435650 90933
rect 434140 90780 434187 90895
rect 435612 90780 435650 90895
rect 434140 90741 435650 90780
rect 509297 90482 509303 90562
rect 509383 90506 510785 90562
rect 509383 90482 509396 90506
rect 434605 89395 435575 89397
rect 434605 89367 436007 89395
rect 434605 89231 434639 89367
rect 435961 89231 436007 89367
rect 434605 89197 436007 89231
rect 509224 88119 509230 88171
rect 509282 88161 509288 88171
rect 509282 88125 510777 88161
rect 509282 88119 509288 88125
rect 509141 85702 509147 85754
rect 509199 85746 509205 85754
rect 509199 85710 510788 85746
rect 509199 85702 509205 85710
rect 430738 83353 444513 83354
rect 430738 83131 444583 83353
rect 427887 82532 428279 82593
rect 427342 81409 427744 81455
rect 427342 80611 427385 81409
rect 427699 80611 427744 81409
rect 427342 80571 427744 80611
rect 427887 80638 427915 82532
rect 428234 80638 428279 82532
rect 427887 80581 428279 80638
rect 435296 81729 436441 82160
rect 444379 82155 444583 83131
rect 435296 80187 435607 81729
rect 439496 81715 441041 82150
rect 444379 81723 445464 82155
rect 439505 81158 440009 81590
rect 444006 81160 444394 81595
rect 445372 81160 445480 81595
rect 439845 78563 440009 81158
rect 385201 78203 385251 78483
rect 385200 78197 385252 78203
rect 389000 78188 389336 78193
rect 398252 78188 398588 78193
rect 402878 78188 403214 78193
rect 407504 78188 407840 78193
rect 412130 78188 412466 78193
rect 416756 78188 417092 78193
rect 421382 78188 421718 78193
rect 426008 78188 426344 78193
rect 430934 78188 431270 78193
rect 435260 78188 435596 78193
rect 385200 78139 385252 78145
rect 435839 77782 435889 78547
rect 439700 78404 440009 78563
rect 444230 78560 444394 81160
rect 448482 81158 449843 81590
rect 440257 78495 440307 78547
rect 440257 78445 440507 78495
rect 435838 77776 435890 77782
rect 435838 77718 435890 77724
rect 374945 74430 375817 74594
rect 374945 73096 375109 74430
rect 439700 70536 439864 78404
rect 440056 78188 440392 78193
rect 440457 77954 440507 78445
rect 444230 78402 444509 78560
rect 444791 78533 444841 78543
rect 444792 78483 445241 78533
rect 440456 77948 440508 77954
rect 440456 77890 440508 77896
rect 444345 70162 444509 78402
rect 444682 78188 445018 78193
rect 445191 78046 445241 78483
rect 449138 78188 449474 78193
rect 445190 78040 445242 78046
rect 445190 77982 445242 77988
rect 449679 74676 449843 81158
rect 507788 80572 508009 84433
rect 551840 84395 551968 95317
rect 552249 94265 556571 94393
rect 559056 94350 560028 95103
rect 552249 84395 552377 94265
rect 563885 94246 564013 95317
rect 567098 94177 568070 94583
rect 568836 88992 568864 89004
rect 568824 88986 568876 88992
rect 568824 88928 568876 88934
rect 509739 83844 510951 83864
rect 509739 83681 509759 83844
rect 510920 83681 510951 83844
rect 509739 83662 510951 83681
rect 509748 82704 510960 82721
rect 509748 82541 509771 82704
rect 510932 82541 510960 82704
rect 509748 82519 510960 82541
rect 550773 82691 551644 82693
rect 550773 82652 551778 82691
rect 550773 82332 550814 82652
rect 551597 82332 551778 82652
rect 550773 82281 551778 82332
rect 515268 80572 515489 81142
rect 526734 80586 526934 81086
rect 536458 80799 536658 81088
rect 536458 80599 537417 80799
rect 546152 80777 546352 81086
rect 507788 80351 515489 80572
rect 507538 79940 507590 79946
rect 507538 79882 507590 79888
rect 507462 79275 507498 79286
rect 507454 79269 507506 79275
rect 507454 79211 507506 79217
rect 507378 79191 507414 79202
rect 507370 79185 507422 79191
rect 507370 79127 507422 79133
rect 507294 79107 507330 79118
rect 507286 79101 507338 79107
rect 507286 79043 507338 79049
rect 507210 79023 507246 79034
rect 507202 79017 507254 79023
rect 507202 78959 507254 78965
rect 507126 78939 507162 78950
rect 448957 74512 449843 74676
rect 448957 74121 449121 74512
rect 289996 62335 290167 69140
rect 290501 62854 290672 69651
rect 292076 61947 292112 61951
rect 292066 61941 292118 61947
rect 292066 61883 292118 61889
rect 289941 61503 289993 61509
rect 289941 61445 289993 61451
rect 289773 61341 289825 61347
rect 289773 61283 289825 61289
rect 289781 5086 289817 61283
rect 289860 61257 289912 61263
rect 289860 61199 289912 61205
rect 289865 5170 289901 61199
rect 289949 5254 289985 61445
rect 290025 61422 290077 61428
rect 290025 61364 290077 61370
rect 290033 5338 290069 61364
rect 292076 19808 292112 61883
rect 292150 61857 292202 61863
rect 292150 61799 292202 61805
rect 292160 20807 292196 61799
rect 292320 61523 292372 61529
rect 292320 61465 292372 61471
rect 292236 61270 292288 61276
rect 292236 61212 292288 61218
rect 292244 21818 292280 61212
rect 292328 22797 292364 61465
rect 292404 61437 292456 61443
rect 292404 61379 292456 61385
rect 292412 23808 292448 61379
rect 292485 61353 292537 61359
rect 292485 61295 292537 61301
rect 292496 24819 292532 61295
rect 319472 60232 319659 67064
rect 320323 60259 320510 67575
rect 340631 61780 340667 61787
rect 340623 61774 340675 61780
rect 340623 61716 340675 61722
rect 340547 61696 340583 61703
rect 340539 61690 340591 61696
rect 340539 61632 340591 61638
rect 340463 61612 340499 61617
rect 340455 61606 340507 61612
rect 340455 61548 340507 61554
rect 320323 60001 320333 60259
rect 340463 26543 340499 61548
rect 339786 26507 340499 26543
rect 340547 25744 340583 61632
rect 339781 25708 340583 25744
rect 340631 24935 340667 61716
rect 339765 24899 340667 24935
rect 341058 61125 341158 61131
rect 292496 24783 292985 24819
rect 292412 23772 293010 23808
rect 292328 22761 293010 22797
rect 292244 21782 292991 21818
rect 292160 20771 293036 20807
rect 292076 19772 293017 19808
rect 294461 19081 295062 19197
rect 294461 16433 294545 19081
rect 295010 16433 295062 19081
rect 341058 17906 341158 61025
rect 342790 59266 342918 62659
rect 342790 56186 342918 58606
rect 343046 56234 343174 62548
rect 343302 59266 343430 63190
rect 343302 56186 343430 58606
rect 343558 56534 343686 63050
rect 343814 59266 343942 63721
rect 343814 56186 343942 58606
rect 344070 56830 344198 63544
rect 344326 59266 344454 64204
rect 344326 56186 344454 58606
rect 344582 57102 344710 64038
rect 344838 59266 344966 64752
rect 344838 56186 344966 58606
rect 345094 57436 345222 64556
rect 345350 59266 345478 65750
rect 345350 56186 345478 58606
rect 345606 57698 345734 65560
rect 345862 59266 345990 65750
rect 345862 56186 345990 58606
rect 346118 57990 346246 64970
rect 346374 59266 346502 69839
rect 346374 56186 346502 58606
rect 346630 58308 346758 69670
rect 346886 59266 347014 69839
rect 347142 58616 347270 69112
rect 347398 59266 347526 69291
rect 346886 56186 347014 58606
rect 347398 56186 347526 58606
rect 348422 59266 348550 66732
rect 348422 56038 348550 58606
rect 348678 57494 348806 66602
rect 348934 59266 349062 66732
rect 348934 56038 349062 58606
rect 349190 57798 349318 66054
rect 349446 59266 349574 67215
rect 349446 56038 349574 58606
rect 349702 58090 349830 67088
rect 349958 59266 350086 67923
rect 349958 56038 350086 58606
rect 350214 58382 350342 67590
rect 350470 59266 350598 68325
rect 350726 58682 350854 68084
rect 350982 59266 351110 68857
rect 350470 56038 350598 58606
rect 351238 58970 351366 68602
rect 351494 59266 351622 68857
rect 350982 56038 351110 58606
rect 351494 56038 351622 58606
rect 352133 59225 354006 59265
rect 352133 58638 352180 59225
rect 353960 58638 354006 59225
rect 352133 58603 354006 58638
rect 364081 58422 364211 68617
rect 364628 58777 364758 68087
rect 385990 63293 386042 63299
rect 385990 63235 386042 63241
rect 374013 62222 374065 62228
rect 374013 62164 374065 62170
rect 354372 54482 354408 54494
rect 354362 54476 354414 54482
rect 354362 54418 354414 54424
rect 354288 49850 354324 49862
rect 354284 49844 354336 49850
rect 354284 49786 354336 49792
rect 353784 45218 353820 45228
rect 353772 45212 353824 45218
rect 353772 45154 353824 45160
rect 353196 42666 353232 42670
rect 353188 42660 353240 42666
rect 353188 42602 353240 42608
rect 353028 37688 353064 37692
rect 353020 37682 353072 37688
rect 353020 37624 353072 37630
rect 352860 32724 352896 32730
rect 352852 32718 352904 32724
rect 352852 32660 352904 32666
rect 352692 27742 352728 27754
rect 352684 27736 352736 27742
rect 352684 27678 352736 27684
rect 352572 18348 352624 18354
rect 352572 18290 352624 18296
rect 341058 17816 341063 17906
rect 341153 17816 341158 17906
rect 341058 17811 341158 17816
rect 341063 17807 341153 17811
rect 352580 17790 352616 18290
rect 352572 17784 352624 17790
rect 352572 17726 352624 17732
rect 352692 17682 352728 27678
rect 352776 27438 352812 27448
rect 352768 27432 352820 27438
rect 352768 27374 352820 27380
rect 352776 17766 352812 27374
rect 352860 17850 352896 32660
rect 352944 32434 352980 32442
rect 352936 32428 352988 32434
rect 352936 32370 352988 32376
rect 352944 17934 352980 32370
rect 353028 18018 353064 37624
rect 353112 37400 353148 37408
rect 353104 37394 353156 37400
rect 353104 37336 353156 37342
rect 353112 18102 353148 37336
rect 353196 18186 353232 42602
rect 353280 42382 353316 42390
rect 353272 42376 353324 42382
rect 353272 42318 353324 42324
rect 353280 18270 353316 42318
rect 353700 39432 353736 39450
rect 353696 39426 353748 39432
rect 353696 39368 353748 39374
rect 353532 22756 353568 22762
rect 353524 22750 353576 22756
rect 353524 22692 353576 22698
rect 353532 18522 353568 22692
rect 353616 22462 353652 22468
rect 353608 22456 353660 22462
rect 353608 22398 353660 22404
rect 353616 18606 353652 22398
rect 353700 18690 353736 39368
rect 353784 18774 353820 45154
rect 353868 34436 353904 34454
rect 353858 34430 353910 34436
rect 353858 34372 353910 34378
rect 353868 18858 353904 34372
rect 353952 29490 353988 29498
rect 353944 29484 353996 29490
rect 353944 29426 353996 29432
rect 353952 18942 353988 29426
rect 354036 24522 354072 24538
rect 354020 24470 354026 24522
rect 354078 24470 354084 24522
rect 354036 19026 354072 24470
rect 354120 19624 354156 19630
rect 354110 19618 354162 19624
rect 354110 19560 354162 19566
rect 354120 19110 354156 19560
rect 354204 19504 354240 19512
rect 354194 19498 354246 19504
rect 354188 19446 354194 19498
rect 354246 19446 354252 19498
rect 354194 19440 354246 19446
rect 354204 19194 354240 19440
rect 354288 19278 354324 49786
rect 354372 19362 354408 54418
rect 374021 48931 374057 62164
rect 374135 62138 374187 62144
rect 374135 62080 374187 62086
rect 374013 48925 374065 48931
rect 374013 48867 374065 48873
rect 374143 48826 374179 62080
rect 374254 61185 374306 61191
rect 374254 61127 374306 61133
rect 374135 48820 374187 48826
rect 374135 48762 374187 48768
rect 374262 48722 374298 61127
rect 374254 48716 374306 48722
rect 374254 48658 374306 48664
rect 385998 44160 386034 63235
rect 391306 61008 391358 61014
rect 391306 60950 391358 60956
rect 385998 44124 386234 44160
rect 385241 43716 386119 43750
rect 385241 43242 385274 43716
rect 386087 43242 386119 43716
rect 385241 43211 386119 43242
rect 386198 42399 386234 44124
rect 385408 42363 386234 42399
rect 384012 41614 385956 41662
rect 384012 41169 384078 41614
rect 385891 41169 385956 41614
rect 384012 41112 385956 41169
rect 367616 40205 367625 40312
rect 367732 40309 367741 40312
rect 367732 40205 367960 40309
rect 391314 40264 391350 60950
rect 385529 40228 391350 40264
rect 391672 45630 392309 45646
rect 367616 40202 367960 40205
rect 384352 39723 385786 39728
rect 391672 39723 392309 45018
rect 392687 44185 392827 60753
rect 405577 60598 405730 61812
rect 407384 61667 407508 69578
rect 405935 61543 407508 61667
rect 405935 60564 406059 61543
rect 411998 61357 412122 69121
rect 453490 64908 453824 78632
rect 454262 78528 454298 78600
rect 454262 78492 454428 78528
rect 454392 77870 454428 78492
rect 454384 77864 454436 77870
rect 454384 77806 454436 77812
rect 458146 74148 458456 78894
rect 458778 78288 458814 78600
rect 458770 78282 458822 78288
rect 458770 78224 458822 78230
rect 458590 78188 458926 78193
rect 462662 73109 462972 78894
rect 467178 78761 467488 78894
rect 463294 78515 463330 78600
rect 463294 78479 463630 78515
rect 463116 78188 463452 78193
rect 463594 77622 463630 78479
rect 467178 78451 467699 78761
rect 467810 78515 467846 78598
rect 467811 78479 468276 78515
rect 463586 77616 463638 77622
rect 463586 77558 463638 77564
rect 467389 68020 467699 78451
rect 467842 78188 468178 78193
rect 468240 77450 468276 78479
rect 471694 78231 472004 78894
rect 471694 77921 472351 78231
rect 472468 78188 472804 78193
rect 468232 77444 468284 77450
rect 468232 77386 468284 77392
rect 472041 66999 472351 77921
rect 476636 65433 476974 78937
rect 507118 78933 507170 78939
rect 481494 78657 481804 78894
rect 477094 78188 477430 78193
rect 477534 77702 477570 78608
rect 481274 78313 481804 78657
rect 482050 78556 482286 78592
rect 477526 77696 477578 77702
rect 477526 77638 477578 77644
rect 481274 74643 481584 78313
rect 481720 78188 482056 78193
rect 482250 78124 482286 78556
rect 482242 78118 482294 78124
rect 482242 78060 482294 78066
rect 485870 73613 486180 78894
rect 486566 78570 486902 78606
rect 486346 78188 486682 78193
rect 486866 77538 486902 78570
rect 486858 77532 486910 77538
rect 486858 77474 486910 77480
rect 490526 68509 490836 78894
rect 491082 78619 491118 78620
rect 491082 78583 491518 78619
rect 490972 78188 491308 78193
rect 491482 77370 491518 78583
rect 491474 77364 491526 77370
rect 491474 77306 491526 77312
rect 495042 67475 495352 78913
rect 507118 78875 507170 78881
rect 507042 78855 507078 78866
rect 507034 78849 507086 78855
rect 507034 78791 507086 78797
rect 506958 78771 506994 78782
rect 506950 78765 507002 78771
rect 506950 78707 507002 78713
rect 506874 78687 506910 78698
rect 506866 78681 506918 78687
rect 506866 78623 506918 78629
rect 495598 78188 495934 78193
rect 499924 78188 500260 78193
rect 506874 68184 506910 78623
rect 506958 68268 506994 78707
rect 507042 68352 507078 78791
rect 507126 68436 507162 78875
rect 507210 68520 507246 78959
rect 507294 68604 507330 79043
rect 507378 68688 507414 79127
rect 507462 68772 507498 79211
rect 507546 68856 507582 79882
rect 507622 79857 507674 79863
rect 507622 79799 507674 79805
rect 507630 68940 507666 79799
rect 507715 79779 507751 79787
rect 507707 79773 507759 79779
rect 507707 79715 507759 79721
rect 507715 69025 507751 79715
rect 507799 79694 507835 79703
rect 507791 79688 507843 79694
rect 507791 79630 507843 79636
rect 507799 69109 507835 79630
rect 507883 79610 507919 79619
rect 507875 79604 507927 79610
rect 507875 79546 507927 79552
rect 507883 69193 507919 79546
rect 507967 79527 508003 79535
rect 507959 79521 508011 79527
rect 507959 79463 508011 79469
rect 507967 69277 508003 79463
rect 508051 79441 508087 79451
rect 508043 79435 508095 79441
rect 508043 79377 508095 79383
rect 508051 69361 508087 79377
rect 508135 79358 508171 79367
rect 508127 79352 508179 79358
rect 537217 79354 537417 80599
rect 551370 80419 551778 82281
rect 556103 82061 556231 82138
rect 555615 81648 556574 82061
rect 563725 82027 563853 82079
rect 555613 81520 556574 81648
rect 555615 81492 556574 81520
rect 559056 81184 560026 82024
rect 563646 81555 564616 82027
rect 567100 80438 568070 82158
rect 543134 80304 544745 80307
rect 543134 80189 548059 80304
rect 543134 79844 543189 80189
rect 544669 79986 548059 80189
rect 544669 79846 544751 79986
rect 568836 79893 568864 88928
rect 568948 88878 568976 88888
rect 568936 88872 568988 88878
rect 568936 88814 568988 88820
rect 566822 79865 568864 79893
rect 544669 79844 544731 79846
rect 543134 79804 544731 79844
rect 508127 79294 508179 79300
rect 508135 69445 508171 79294
rect 510410 78460 510446 78466
rect 510402 78454 510454 78460
rect 510402 78396 510454 78402
rect 510326 78376 510362 78382
rect 510318 78370 510370 78376
rect 510318 78312 510370 78318
rect 510242 78292 510278 78298
rect 510234 78286 510286 78292
rect 510234 78228 510286 78234
rect 510158 78208 510194 78214
rect 510150 78202 510202 78208
rect 510150 78144 510202 78150
rect 510074 78124 510110 78130
rect 510066 78118 510118 78124
rect 510066 78060 510118 78066
rect 509990 78040 510026 78046
rect 509982 78034 510034 78040
rect 509982 77976 510034 77982
rect 509906 77956 509942 77962
rect 509898 77950 509950 77956
rect 509898 77892 509950 77898
rect 509822 77872 509858 77878
rect 509814 77866 509866 77872
rect 509814 77808 509866 77814
rect 509738 77788 509774 77794
rect 509730 77782 509782 77788
rect 509730 77724 509782 77730
rect 509654 77704 509690 77710
rect 509646 77698 509698 77704
rect 509646 77640 509698 77646
rect 509570 77620 509606 77626
rect 509562 77614 509614 77620
rect 509562 77556 509614 77562
rect 509486 77536 509522 77542
rect 509478 77530 509530 77536
rect 509478 77472 509530 77478
rect 509402 77452 509438 77458
rect 509394 77446 509446 77452
rect 509394 77388 509446 77394
rect 509318 77368 509354 77374
rect 509310 77362 509362 77368
rect 509310 77304 509362 77310
rect 509318 69548 509354 77304
rect 509402 69632 509438 77388
rect 509486 69716 509522 77472
rect 509570 69800 509606 77556
rect 509654 69884 509690 77640
rect 509738 69968 509774 77724
rect 509822 70052 509858 77808
rect 509906 70136 509942 77892
rect 509990 70220 510026 77976
rect 510074 70304 510110 78060
rect 510158 70388 510194 78144
rect 510242 70472 510278 78228
rect 510326 70556 510362 78312
rect 510410 70640 510446 78396
rect 528478 78316 528514 78333
rect 528470 78310 528522 78316
rect 528470 78252 528522 78258
rect 528394 78232 528430 78249
rect 528386 78226 528438 78232
rect 528386 78168 528438 78174
rect 528310 78148 528346 78165
rect 528302 78142 528354 78148
rect 528302 78084 528354 78090
rect 528226 78064 528262 78081
rect 528218 78058 528270 78064
rect 528218 78000 528270 78006
rect 528142 77980 528178 77997
rect 528134 77974 528186 77980
rect 528134 77916 528186 77922
rect 528058 77896 528094 77913
rect 528050 77890 528102 77896
rect 528050 77832 528102 77838
rect 527974 77812 528010 77829
rect 527966 77806 528018 77812
rect 527966 77748 528018 77754
rect 527890 77728 527926 77745
rect 527882 77722 527934 77728
rect 527882 77664 527934 77670
rect 527806 77644 527842 77661
rect 527798 77638 527850 77644
rect 527798 77580 527850 77586
rect 527722 77560 527758 77577
rect 527714 77554 527766 77560
rect 527714 77496 527766 77502
rect 527422 77198 527458 77206
rect 527414 77192 527466 77198
rect 527414 77134 527466 77140
rect 526846 77114 526882 77120
rect 526838 77108 526890 77114
rect 526838 77050 526890 77056
rect 526486 77030 526522 77032
rect 526478 77024 526530 77030
rect 526478 76966 526530 76972
rect 525334 76948 525370 76962
rect 525326 76942 525378 76948
rect 525326 76884 525378 76890
rect 525262 76274 525298 76280
rect 525254 76268 525306 76274
rect 525254 76210 525306 76216
rect 524830 75854 524866 75862
rect 524822 75848 524874 75854
rect 524822 75790 524874 75796
rect 510410 70604 523546 70640
rect 510326 70520 523462 70556
rect 510242 70436 523378 70472
rect 510158 70352 523294 70388
rect 510074 70268 523210 70304
rect 509990 70184 523126 70220
rect 509906 70100 523042 70136
rect 509822 70016 522958 70052
rect 509738 69932 522874 69968
rect 509654 69848 522790 69884
rect 509570 69764 522706 69800
rect 509486 69680 522622 69716
rect 509402 69596 522538 69632
rect 509318 69512 522454 69548
rect 508135 69409 522071 69445
rect 508051 69325 521987 69361
rect 507967 69241 521903 69277
rect 507883 69157 521819 69193
rect 507799 69073 521735 69109
rect 507715 68989 521651 69025
rect 507630 68904 521566 68940
rect 507546 68820 521482 68856
rect 507462 68736 521398 68772
rect 507378 68652 521314 68688
rect 507294 68568 521230 68604
rect 507210 68484 521146 68520
rect 507126 68400 521062 68436
rect 507042 68316 520978 68352
rect 506958 68232 520894 68268
rect 506874 68148 520810 68184
rect 416050 63216 416086 63219
rect 416042 63210 416094 63216
rect 480559 63214 480595 63226
rect 416042 63152 416094 63158
rect 480551 63208 480603 63214
rect 415966 63132 416002 63142
rect 415958 63126 416010 63132
rect 415958 63068 416010 63074
rect 415882 63048 415918 63057
rect 415874 63042 415926 63048
rect 415874 62984 415926 62990
rect 415798 62963 415834 62968
rect 415790 62957 415842 62963
rect 415790 62899 415842 62905
rect 415714 61870 415750 61874
rect 415706 61864 415758 61870
rect 415706 61806 415758 61812
rect 406245 61233 412122 61357
rect 406245 60588 406369 61233
rect 406677 59916 407807 59944
rect 406677 59616 406725 59916
rect 407761 59616 407807 59916
rect 406677 59583 407807 59616
rect 401933 45507 401969 46594
rect 402220 45614 402256 46470
rect 403880 46464 404079 46486
rect 403880 46006 403905 46464
rect 404057 46006 404079 46464
rect 403880 45980 404079 46006
rect 404186 46458 404385 46486
rect 404186 46000 404206 46458
rect 404358 46000 404385 46458
rect 404186 45980 404385 46000
rect 415714 45902 415750 61806
rect 415706 45896 415758 45902
rect 415706 45838 415758 45844
rect 415714 45834 415750 45838
rect 415798 45811 415834 62899
rect 415790 45805 415842 45811
rect 415790 45747 415842 45753
rect 415798 45741 415834 45747
rect 415882 45725 415918 62984
rect 415874 45719 415926 45725
rect 415874 45661 415926 45667
rect 415882 45652 415918 45661
rect 415966 45627 416002 63068
rect 402900 45614 402906 45622
rect 402220 45578 402906 45614
rect 402900 45570 402906 45578
rect 402958 45570 402964 45622
rect 415958 45621 416010 45627
rect 415958 45563 416010 45569
rect 415966 45558 416002 45563
rect 416050 45520 416086 63152
rect 480551 63150 480603 63156
rect 421035 51919 421805 51943
rect 421035 51916 421070 51919
rect 420956 51773 421070 51916
rect 421767 51773 421805 51919
rect 420956 51748 421805 51773
rect 421035 51738 421805 51748
rect 422027 51471 422210 61869
rect 430608 61622 431282 61628
rect 429754 61588 430580 61590
rect 429754 61522 429774 61588
rect 430184 61522 430580 61588
rect 429754 61518 430580 61522
rect 422513 60346 422565 60352
rect 422513 60288 422565 60294
rect 422521 60269 422558 60288
rect 420904 51288 422210 51471
rect 416981 49325 417583 49462
rect 402902 45507 402908 45515
rect 401933 45471 402908 45507
rect 402902 45463 402908 45471
rect 402960 45463 402966 45515
rect 416042 45514 416094 45520
rect 416042 45456 416094 45462
rect 416050 45451 416086 45456
rect 416981 44430 417118 49325
rect 421021 48814 422062 48919
rect 420994 48487 421764 48507
rect 420994 48341 421046 48487
rect 421743 48341 421764 48487
rect 420994 48317 421764 48341
rect 420754 47158 421778 47190
rect 420754 47148 421781 47158
rect 420754 47023 420803 47148
rect 421743 47023 421781 47148
rect 420754 46988 421781 47023
rect 420747 46173 421736 46211
rect 420747 46034 420789 46173
rect 421670 46034 421736 46173
rect 420747 46003 421736 46034
rect 421950 44616 422062 48814
rect 422522 47576 422558 60269
rect 422514 47570 422566 47576
rect 422514 47512 422566 47518
rect 384352 39680 392309 39723
rect 384352 39126 384400 39680
rect 385734 39126 392309 39680
rect 384352 39086 392309 39126
rect 384352 39078 385786 39086
rect 430508 37750 430580 61518
rect 430094 37678 430580 37750
rect 430608 61564 430758 61622
rect 431270 61564 431282 61622
rect 430608 61560 431282 61564
rect 430608 36998 430676 61560
rect 430717 61522 430769 61528
rect 430717 61464 430769 61470
rect 430084 36930 430676 36998
rect 393739 32731 395092 32753
rect 393739 32474 393779 32731
rect 394848 32474 395092 32731
rect 430724 32645 430760 61464
rect 430808 61444 430844 61447
rect 430800 61438 430852 61444
rect 430800 61380 430852 61386
rect 430265 32609 430760 32645
rect 393739 32443 395092 32474
rect 430255 31890 430749 31916
rect 430715 31573 430749 31890
rect 430255 31541 430749 31573
rect 430808 31107 430844 61380
rect 446720 45172 446789 45187
rect 436476 44757 436556 45046
rect 446720 44680 446789 44838
rect 446772 44628 446789 44680
rect 446720 44619 446789 44628
rect 446880 45172 446949 45187
rect 446880 44512 446949 44838
rect 446880 44460 446884 44512
rect 446936 44460 446949 44512
rect 446880 44453 446949 44460
rect 447040 45172 447109 45187
rect 447040 44344 447109 44838
rect 447040 44292 447043 44344
rect 447095 44292 447109 44344
rect 447040 44273 447109 44292
rect 447200 45172 447269 45187
rect 447200 44176 447269 44838
rect 447200 44124 447207 44176
rect 447259 44124 447269 44176
rect 447200 44113 447269 44124
rect 447360 45172 447429 45187
rect 447360 44008 447429 44838
rect 447360 43956 447365 44008
rect 447417 43956 447429 44008
rect 447360 43949 447429 43956
rect 447520 45172 447589 45187
rect 447520 43840 447589 44838
rect 447520 43788 447524 43840
rect 447576 43788 447589 43840
rect 447520 43774 447589 43788
rect 447680 45172 447749 45187
rect 447680 43672 447749 44838
rect 447680 43620 447688 43672
rect 447740 43620 447749 43672
rect 447680 43607 447749 43620
rect 447840 45172 447909 45187
rect 447840 43504 447909 44838
rect 451596 45175 451665 45190
rect 451596 43588 451665 44841
rect 451756 45175 451825 45190
rect 451756 43756 451825 44841
rect 451916 45175 451985 45190
rect 451916 43924 451985 44841
rect 452076 45175 452145 45190
rect 452076 44092 452145 44841
rect 452236 45175 452305 45190
rect 452236 44260 452305 44841
rect 452396 45175 452465 45190
rect 452396 44428 452465 44841
rect 452556 45175 452625 45190
rect 452556 44596 452625 44841
rect 452716 45175 452785 45190
rect 452716 44764 452785 44841
rect 480559 44767 480595 63150
rect 480643 63130 480679 63151
rect 480635 63124 480687 63130
rect 480635 63066 480687 63072
rect 452716 44712 452727 44764
rect 452779 44712 452785 44764
rect 452716 44697 452785 44712
rect 480551 44761 480603 44767
rect 480551 44703 480603 44709
rect 480559 44701 480595 44703
rect 480643 44683 480679 63066
rect 480727 63046 480763 63067
rect 480719 63040 480771 63046
rect 480719 62982 480771 62988
rect 480635 44677 480687 44683
rect 480635 44619 480687 44625
rect 480643 44617 480679 44619
rect 480727 44599 480763 62982
rect 480811 62962 480847 62983
rect 480803 62956 480855 62962
rect 480803 62898 480855 62904
rect 452556 44544 452565 44596
rect 452617 44544 452625 44596
rect 452556 44532 452625 44544
rect 480719 44593 480771 44599
rect 480719 44535 480771 44541
rect 480727 44533 480763 44535
rect 480811 44515 480847 62898
rect 480895 62878 480931 62899
rect 480887 62872 480939 62878
rect 480887 62814 480939 62820
rect 480803 44509 480855 44515
rect 480803 44451 480855 44457
rect 480811 44449 480847 44451
rect 480895 44431 480931 62814
rect 480979 62794 481015 62815
rect 480971 62788 481023 62794
rect 480971 62730 481023 62736
rect 452396 44376 452405 44428
rect 452457 44376 452465 44428
rect 452396 44366 452465 44376
rect 480887 44425 480939 44431
rect 480887 44367 480939 44373
rect 480895 44365 480931 44367
rect 480979 44347 481015 62730
rect 481063 62710 481099 62731
rect 481055 62704 481107 62710
rect 481055 62646 481107 62652
rect 480971 44341 481023 44347
rect 480971 44283 481023 44289
rect 480979 44281 481015 44283
rect 481063 44263 481099 62646
rect 481147 62626 481183 62647
rect 481139 62620 481191 62626
rect 481139 62562 481191 62568
rect 452236 44208 452243 44260
rect 452295 44208 452305 44260
rect 452236 44190 452305 44208
rect 481055 44257 481107 44263
rect 481055 44199 481107 44205
rect 481063 44197 481099 44199
rect 481147 44179 481183 62562
rect 481231 62542 481267 62563
rect 481223 62536 481275 62542
rect 481223 62478 481275 62484
rect 485638 62540 519124 62576
rect 481139 44173 481191 44179
rect 481139 44115 481191 44121
rect 481147 44113 481183 44115
rect 481231 44095 481267 62478
rect 481315 62458 481351 62479
rect 481307 62452 481359 62458
rect 481307 62394 481359 62400
rect 452076 44040 452088 44092
rect 452140 44040 452145 44092
rect 452076 44028 452145 44040
rect 481223 44089 481275 44095
rect 481223 44031 481275 44037
rect 481231 44029 481267 44031
rect 481315 44011 481351 62394
rect 481399 62374 481435 62395
rect 481391 62368 481443 62374
rect 481391 62310 481443 62316
rect 481307 44005 481359 44011
rect 481307 43947 481359 43953
rect 481315 43945 481351 43947
rect 481399 43927 481435 62310
rect 481483 62290 481519 62311
rect 481475 62284 481527 62290
rect 481475 62226 481527 62232
rect 451916 43872 451920 43924
rect 451972 43872 451985 43924
rect 451916 43864 451985 43872
rect 481391 43921 481443 43927
rect 481391 43863 481443 43869
rect 481399 43861 481435 43863
rect 481483 43843 481519 62226
rect 481567 62206 481603 62227
rect 481559 62200 481611 62206
rect 481559 62142 481611 62148
rect 481475 43837 481527 43843
rect 481475 43779 481527 43785
rect 481483 43777 481519 43779
rect 481567 43759 481603 62142
rect 481651 62122 481687 62143
rect 481643 62116 481695 62122
rect 481643 62058 481695 62064
rect 451756 43704 451765 43756
rect 451817 43704 451825 43756
rect 451756 43691 451825 43704
rect 481559 43753 481611 43759
rect 481559 43695 481611 43701
rect 481567 43693 481603 43695
rect 481651 43675 481687 62058
rect 481735 62038 481771 62059
rect 481727 62032 481779 62038
rect 481727 61974 481779 61980
rect 481643 43669 481695 43675
rect 481643 43611 481695 43617
rect 481651 43609 481687 43611
rect 481735 43591 481771 61974
rect 481819 61954 481855 61975
rect 481811 61948 481863 61954
rect 481811 61890 481863 61896
rect 451596 43536 451603 43588
rect 451655 43536 451665 43588
rect 451596 43519 451665 43536
rect 481727 43585 481779 43591
rect 481727 43527 481779 43533
rect 481735 43525 481771 43527
rect 481819 43507 481855 61890
rect 481937 60599 481989 60605
rect 481937 60541 481989 60547
rect 447840 43452 447846 43504
rect 447898 43452 447909 43504
rect 447840 43439 447909 43452
rect 481811 43501 481863 43507
rect 481811 43443 481863 43449
rect 481819 43442 481855 43443
rect 451969 42875 459639 43075
rect 451969 41808 452125 42875
rect 459416 41808 459639 42875
rect 451969 41608 459639 41808
rect 472888 42852 480558 43008
rect 472888 41785 473111 42852
rect 480402 41785 480558 42852
rect 472888 41541 480558 41785
rect 481945 36094 481981 60541
rect 482109 44396 482416 44405
rect 482109 44280 482416 44289
rect 478145 36058 481981 36094
rect 482126 31443 482188 44280
rect 483618 44250 483763 61832
rect 485638 61024 485674 62540
rect 485722 62456 519040 62492
rect 485628 61018 485680 61024
rect 485628 60960 485680 60966
rect 485722 60940 485758 62456
rect 485806 62372 518956 62408
rect 485712 60934 485764 60940
rect 485712 60876 485764 60882
rect 485722 60872 485758 60876
rect 485806 60856 485842 62372
rect 485890 62288 518872 62324
rect 485794 60850 485846 60856
rect 485794 60792 485846 60798
rect 485806 60786 485842 60792
rect 485890 60772 485926 62288
rect 485974 62204 518788 62240
rect 485882 60766 485934 60772
rect 485882 60708 485934 60714
rect 485890 60702 485926 60708
rect 485974 60688 486010 62204
rect 486058 62120 518704 62156
rect 485968 60682 486020 60688
rect 485968 60624 486020 60630
rect 485974 60612 486010 60624
rect 486058 60604 486094 62120
rect 486142 62036 518620 62072
rect 486046 60598 486098 60604
rect 486046 60540 486098 60546
rect 486058 60532 486094 60540
rect 486142 60520 486178 62036
rect 486226 61952 518536 61988
rect 486136 60514 486188 60520
rect 486136 60456 486188 60462
rect 486142 60448 486178 60456
rect 486226 60436 486262 61952
rect 486310 61868 518452 61904
rect 486216 60430 486268 60436
rect 486216 60372 486268 60378
rect 486226 60368 486262 60372
rect 486310 60352 486346 61868
rect 486394 61784 518368 61820
rect 486298 60346 486350 60352
rect 486298 60288 486350 60294
rect 486310 60282 486346 60288
rect 486394 60268 486430 61784
rect 486478 61700 518284 61736
rect 486382 60262 486434 60268
rect 486382 60204 486434 60210
rect 486394 60196 486430 60204
rect 486478 60184 486514 61700
rect 518248 60184 518284 61700
rect 518332 60268 518368 61784
rect 518416 60352 518452 61868
rect 518500 60436 518536 61952
rect 518584 60520 518620 62036
rect 518668 60604 518704 62120
rect 518752 60688 518788 62204
rect 518836 60772 518872 62288
rect 518920 60856 518956 62372
rect 519004 60940 519040 62456
rect 519088 61024 519124 62540
rect 519080 61018 519132 61024
rect 519080 60960 519132 60966
rect 519088 60950 519124 60960
rect 518996 60934 519048 60940
rect 518996 60876 519048 60882
rect 519004 60874 519040 60876
rect 518912 60850 518964 60856
rect 518912 60792 518964 60798
rect 518920 60788 518956 60792
rect 518828 60766 518880 60772
rect 518828 60708 518880 60714
rect 518836 60706 518872 60708
rect 518744 60682 518796 60688
rect 518744 60624 518796 60630
rect 518752 60618 518788 60624
rect 518660 60598 518712 60604
rect 518660 60540 518712 60546
rect 518668 60538 518704 60540
rect 518576 60514 518628 60520
rect 518576 60456 518628 60462
rect 518584 60450 518620 60456
rect 518492 60430 518544 60436
rect 518492 60372 518544 60378
rect 518500 60368 518536 60372
rect 518408 60346 518460 60352
rect 518408 60288 518460 60294
rect 518416 60282 518452 60288
rect 518324 60262 518376 60268
rect 518324 60204 518376 60210
rect 518332 60198 518368 60204
rect 486468 60178 486520 60184
rect 486468 60120 486520 60126
rect 518240 60178 518292 60184
rect 518240 60120 518292 60126
rect 478191 31381 482188 31443
rect 430267 31071 430844 31107
rect 392020 29084 394378 29116
rect 392020 28615 392065 29084
rect 392969 28615 394378 29084
rect 392020 28577 394378 28615
rect 520774 25879 520810 68148
rect 520858 25963 520894 68232
rect 520942 26047 520978 68316
rect 521026 26131 521062 68400
rect 521110 26215 521146 68484
rect 521194 26299 521230 68568
rect 521278 26383 521314 68652
rect 521362 26467 521398 68736
rect 521446 26551 521482 68820
rect 521530 26635 521566 68904
rect 521615 26719 521651 68989
rect 521699 26803 521735 69073
rect 521783 26887 521819 69157
rect 521867 26971 521903 69241
rect 521951 27055 521987 69325
rect 522035 27139 522071 69409
rect 522327 61613 522363 61617
rect 522319 61607 522371 61613
rect 522223 61529 522259 61535
rect 522215 61523 522267 61529
rect 522215 61465 522267 61471
rect 522139 61444 522175 61448
rect 522131 61438 522183 61444
rect 522131 61380 522183 61386
rect 522139 49751 522175 61380
rect 522223 49836 522259 61465
rect 522307 61395 522319 61426
rect 522307 61389 522371 61395
rect 522307 50120 522363 61389
rect 522299 50114 522363 50120
rect 522351 49862 522363 50114
rect 522299 49858 522363 49862
rect 522299 49856 522351 49858
rect 522215 49830 522267 49836
rect 522215 49772 522267 49778
rect 522131 49745 522183 49751
rect 522131 49687 522183 49693
rect 522418 36418 522454 69512
rect 522502 36502 522538 69596
rect 522586 36586 522622 69680
rect 522670 36670 522706 69764
rect 522754 36754 522790 69848
rect 522838 36838 522874 69932
rect 522922 36922 522958 70016
rect 523006 37006 523042 70100
rect 523090 37090 523126 70184
rect 523174 37174 523210 70268
rect 523258 37258 523294 70352
rect 523342 37342 523378 70436
rect 523426 37426 523462 70520
rect 523510 37510 523546 70604
rect 524182 65832 524218 65836
rect 524174 65826 524226 65832
rect 524174 65768 524226 65774
rect 523678 65748 523714 65760
rect 523670 65742 523722 65748
rect 523670 65684 523722 65690
rect 523678 40158 523714 65684
rect 523966 65496 524002 65504
rect 523958 65490 524010 65496
rect 523958 65432 524010 65438
rect 523750 65162 523786 65166
rect 523742 65156 523794 65162
rect 523742 65098 523794 65104
rect 523750 40230 523786 65098
rect 523822 64320 523858 64338
rect 523814 64314 523866 64320
rect 523814 64256 523866 64262
rect 523822 40302 523858 64256
rect 523894 63480 523930 63488
rect 523886 63474 523938 63480
rect 523886 63416 523938 63422
rect 523894 40374 523930 63416
rect 523966 40446 524002 65432
rect 524038 64740 524074 64744
rect 524030 64734 524082 64740
rect 524030 64676 524082 64682
rect 524038 40518 524074 64676
rect 524110 63900 524146 63912
rect 524102 63894 524154 63900
rect 524102 63836 524154 63842
rect 524110 40590 524146 63836
rect 524182 40662 524218 65768
rect 524470 65580 524506 65584
rect 524462 65574 524514 65580
rect 524462 65516 524514 65522
rect 524254 65244 524290 65248
rect 524246 65238 524298 65244
rect 524246 65180 524298 65186
rect 524254 40734 524290 65180
rect 524326 64404 524362 64418
rect 524318 64398 524370 64404
rect 524318 64340 524370 64346
rect 524326 40806 524362 64340
rect 524398 63564 524434 63570
rect 524390 63558 524442 63564
rect 524390 63500 524442 63506
rect 524398 40878 524434 63500
rect 524470 40950 524506 65516
rect 524686 64908 524722 64912
rect 524678 64902 524730 64908
rect 524678 64844 524730 64850
rect 524542 64826 524578 64832
rect 524534 64820 524586 64826
rect 524534 64762 524586 64768
rect 524542 41022 524578 64762
rect 524614 63984 524650 63990
rect 524606 63978 524658 63984
rect 524606 63920 524658 63926
rect 524614 41094 524650 63920
rect 524686 41166 524722 64844
rect 524758 64068 524794 64074
rect 524750 64062 524802 64068
rect 524750 64004 524802 64010
rect 524758 41238 524794 64004
rect 524830 41310 524866 75790
rect 525046 75770 525082 75772
rect 525038 75764 525090 75770
rect 525038 75706 525090 75712
rect 524902 64490 524938 64508
rect 524894 64484 524946 64490
rect 524894 64426 524946 64432
rect 524902 41382 524938 64426
rect 524974 63648 525010 63658
rect 524966 63642 525018 63648
rect 524966 63584 525018 63590
rect 524974 41454 525010 63584
rect 525046 41526 525082 75706
rect 525118 64572 525154 64580
rect 525110 64566 525162 64572
rect 525110 64508 525162 64514
rect 525118 41598 525154 64508
rect 525190 63732 525226 63740
rect 525182 63726 525234 63732
rect 525182 63668 525234 63674
rect 525190 41670 525226 63668
rect 525262 41742 525298 76210
rect 525334 41814 525370 76884
rect 525766 76610 525802 76616
rect 525758 76604 525810 76610
rect 525758 76546 525810 76552
rect 525694 75940 525730 75946
rect 525686 75934 525738 75940
rect 525686 75876 525738 75882
rect 525622 75602 525658 75612
rect 525614 75596 525666 75602
rect 525614 75538 525666 75544
rect 525406 75434 525442 75446
rect 525398 75428 525450 75434
rect 525398 75370 525450 75376
rect 525406 41886 525442 75370
rect 525478 64992 525514 64998
rect 525470 64986 525522 64992
rect 525470 64928 525522 64934
rect 525478 41958 525514 64928
rect 525550 64152 525586 64156
rect 525542 64146 525594 64152
rect 525542 64088 525594 64094
rect 525550 42030 525586 64088
rect 525622 42102 525658 75538
rect 525694 42174 525730 75876
rect 525766 42246 525802 76546
rect 526414 76358 526450 76368
rect 526406 76352 526458 76358
rect 526406 76294 526458 76300
rect 526342 75686 526378 75692
rect 526334 75680 526386 75686
rect 526334 75622 526386 75628
rect 525838 65664 525874 65670
rect 525830 65658 525882 65664
rect 525830 65600 525882 65606
rect 525838 42318 525874 65600
rect 526126 65416 526162 65420
rect 526118 65410 526170 65416
rect 526118 65352 526170 65358
rect 525910 65078 525946 65082
rect 525902 65072 525954 65078
rect 525902 65014 525954 65020
rect 525910 42390 525946 65014
rect 525982 64236 526018 64242
rect 525974 64230 526026 64236
rect 525974 64172 526026 64178
rect 525982 42462 526018 64172
rect 526054 63396 526090 63400
rect 526046 63390 526098 63396
rect 526046 63332 526098 63338
rect 526054 42534 526090 63332
rect 526126 42606 526162 65352
rect 526198 64656 526234 64664
rect 526190 64650 526242 64656
rect 526190 64592 526242 64598
rect 526198 42678 526234 64592
rect 526270 63816 526306 63826
rect 526262 63810 526314 63816
rect 526262 63752 526314 63758
rect 526270 42750 526306 63752
rect 526342 42822 526378 75622
rect 526414 42894 526450 76294
rect 526486 42966 526522 76966
rect 526702 76694 526738 76700
rect 526694 76688 526746 76694
rect 526694 76630 526746 76636
rect 526630 76022 526666 76028
rect 526622 76016 526674 76022
rect 526622 75958 526674 75964
rect 526558 75348 526594 75354
rect 526550 75342 526602 75348
rect 526550 75284 526602 75290
rect 526558 43038 526594 75284
rect 526630 43110 526666 75958
rect 526702 43182 526738 76630
rect 526774 76442 526810 76452
rect 526766 76436 526818 76442
rect 526766 76378 526818 76384
rect 526774 43254 526810 76378
rect 526846 43326 526882 77050
rect 527198 76856 527250 76862
rect 527198 76798 527250 76804
rect 527062 76778 527098 76782
rect 527054 76772 527106 76778
rect 527054 76714 527106 76720
rect 526990 76106 527026 76112
rect 526982 76100 527034 76106
rect 526982 76042 527034 76048
rect 526918 75520 526954 75528
rect 526910 75514 526962 75520
rect 526910 75456 526962 75462
rect 526918 43398 526954 75456
rect 526990 43470 527026 76042
rect 527062 43542 527098 76714
rect 527134 76192 527170 76198
rect 527126 76186 527178 76192
rect 527126 76128 527178 76134
rect 527134 43614 527170 76128
rect 527206 43686 527242 76798
rect 527350 76526 527386 76530
rect 527342 76520 527394 76526
rect 527342 76462 527394 76468
rect 527278 65328 527314 65332
rect 527270 65322 527322 65328
rect 527270 65264 527322 65270
rect 527278 43758 527314 65264
rect 527350 43830 527386 76462
rect 527422 43902 527458 77134
rect 527722 44904 527758 77496
rect 527806 44988 527842 77580
rect 527890 45072 527926 77664
rect 527974 45156 528010 77748
rect 528058 45240 528094 77832
rect 528142 45324 528178 77916
rect 528226 45408 528262 78000
rect 528310 45492 528346 78084
rect 528394 45576 528430 78168
rect 528478 45660 528514 78252
rect 528646 77381 528682 77395
rect 528638 77375 528690 77381
rect 528638 77317 528690 77323
rect 528562 77285 528598 77286
rect 528557 77279 528609 77285
rect 528557 77221 528609 77227
rect 528562 45744 528598 77221
rect 528646 45828 528682 77317
rect 546101 75164 546229 78655
rect 546577 75662 546705 78691
rect 547058 74676 547186 78320
rect 547551 74207 547679 77595
rect 544438 63298 544474 63311
rect 544430 63292 544482 63298
rect 544430 63234 544482 63240
rect 544354 63214 544390 63227
rect 544346 63208 544398 63214
rect 544346 63150 544398 63156
rect 544270 63130 544306 63143
rect 544262 63124 544314 63130
rect 544262 63066 544314 63072
rect 544186 63046 544222 63059
rect 544178 63040 544230 63046
rect 544178 62982 544230 62988
rect 544102 62962 544138 62975
rect 544094 62956 544146 62962
rect 544094 62898 544146 62904
rect 544018 62878 544054 62891
rect 544010 62872 544062 62878
rect 544010 62814 544062 62820
rect 543934 62794 543970 62807
rect 543926 62788 543978 62794
rect 543926 62730 543978 62736
rect 543850 62710 543886 62723
rect 543842 62704 543894 62710
rect 543842 62646 543894 62652
rect 543766 62626 543802 62639
rect 543758 62620 543810 62626
rect 543758 62562 543810 62568
rect 543682 62542 543718 62555
rect 543674 62536 543726 62542
rect 543674 62478 543726 62484
rect 543598 62458 543634 62471
rect 543590 62452 543642 62458
rect 543590 62394 543642 62400
rect 543514 62374 543550 62387
rect 543506 62368 543558 62374
rect 543506 62310 543558 62316
rect 543430 62290 543466 62303
rect 543422 62284 543474 62290
rect 543422 62226 543474 62232
rect 543346 62206 543382 62219
rect 543338 62200 543390 62206
rect 543338 62142 543390 62148
rect 543262 62122 543298 62135
rect 543254 62116 543306 62122
rect 543254 62058 543306 62064
rect 543178 62038 543214 62051
rect 543170 62032 543222 62038
rect 543170 61974 543222 61980
rect 543094 61954 543130 61967
rect 543086 61948 543138 61954
rect 543086 61890 543138 61896
rect 543010 61870 543046 61883
rect 543002 61864 543054 61870
rect 543002 61806 543054 61812
rect 542926 61786 542962 61799
rect 542918 61780 542970 61786
rect 542918 61722 542970 61728
rect 542842 61702 542878 61715
rect 542834 61696 542886 61702
rect 542834 61638 542886 61644
rect 542750 61354 542802 61360
rect 542750 61296 542802 61302
rect 542674 61276 542710 61289
rect 542666 61270 542718 61276
rect 542666 61212 542718 61218
rect 542590 61192 542626 61205
rect 542582 61186 542634 61192
rect 542582 61128 542634 61134
rect 542506 61108 542542 61121
rect 542498 61102 542550 61108
rect 542498 61044 542550 61050
rect 542422 61024 542458 61037
rect 542414 61018 542466 61024
rect 542414 60960 542466 60966
rect 542338 60940 542374 60953
rect 542330 60934 542382 60940
rect 542330 60876 542382 60882
rect 542254 60856 542290 60869
rect 542246 60850 542298 60856
rect 542246 60792 542298 60798
rect 542170 60772 542206 60785
rect 542162 60766 542214 60772
rect 542162 60708 542214 60714
rect 542086 60688 542122 60701
rect 542078 60682 542130 60688
rect 542078 60624 542130 60630
rect 542002 60604 542038 60617
rect 541994 60598 542046 60604
rect 541994 60540 542046 60546
rect 541918 60520 541954 60533
rect 541910 60514 541962 60520
rect 541910 60456 541962 60462
rect 541834 60436 541870 60449
rect 541826 60430 541878 60436
rect 541826 60372 541878 60378
rect 541750 60352 541786 60365
rect 541742 60346 541794 60352
rect 541742 60288 541794 60294
rect 541666 60268 541702 60281
rect 541658 60262 541710 60268
rect 541658 60204 541710 60210
rect 541582 60184 541618 60197
rect 541574 60178 541626 60184
rect 541574 60120 541626 60126
rect 541582 56507 541618 60120
rect 541666 56591 541702 60204
rect 541750 56675 541786 60288
rect 541834 56759 541870 60372
rect 541918 56843 541954 60456
rect 542002 56927 542038 60540
rect 542086 57011 542122 60624
rect 542170 57095 542206 60708
rect 542254 57179 542290 60792
rect 542338 57263 542374 60876
rect 542422 57347 542458 60960
rect 542506 57431 542542 61044
rect 542590 57515 542626 61128
rect 542674 57599 542710 61212
rect 542758 57683 542794 61296
rect 542842 57767 542878 61638
rect 542926 57851 542962 61722
rect 543010 57935 543046 61806
rect 543094 58019 543130 61890
rect 543178 58103 543214 61974
rect 543262 58187 543298 62058
rect 543346 58271 543382 62142
rect 543430 58355 543466 62226
rect 543514 58439 543550 62310
rect 543598 58523 543634 62394
rect 543682 58607 543718 62478
rect 543766 58691 543802 62562
rect 543850 58775 543886 62646
rect 543934 58859 543970 62730
rect 544018 58943 544054 62814
rect 544102 59027 544138 62898
rect 544186 59111 544222 62982
rect 544270 59195 544306 63066
rect 544354 59279 544390 63150
rect 544438 59363 544474 63234
rect 551206 60908 551870 61112
rect 550995 60849 551870 60908
rect 547846 60451 547882 60500
rect 547246 60415 547882 60451
rect 547246 60374 547282 60415
rect 547918 60382 547954 60497
rect 547318 60346 547954 60382
rect 547318 60256 547354 60346
rect 547990 60310 548026 60495
rect 547390 60274 548026 60310
rect 547390 60138 547426 60274
rect 548062 60237 548098 60495
rect 547462 60202 548098 60237
rect 550881 60476 551870 60849
rect 562697 60665 564300 60715
rect 550881 60475 552176 60476
rect 547462 60201 548096 60202
rect 547462 60016 547498 60201
rect 550881 60069 552178 60475
rect 550881 59817 552176 60069
rect 552478 59724 552514 60508
rect 552550 59836 552586 60496
rect 552622 59926 552658 60512
rect 552694 60036 552730 60510
rect 555796 60044 556768 60324
rect 557110 60116 557146 60547
rect 557182 60228 557218 60547
rect 557254 60342 557290 60547
rect 557326 60452 557362 60547
rect 561020 60518 561048 60540
rect 561010 60512 561062 60518
rect 561010 60454 561062 60460
rect 559248 59964 560220 60064
rect 544438 59327 544928 59363
rect 544354 59243 544844 59279
rect 544270 59159 544760 59195
rect 544186 59075 544676 59111
rect 544102 58991 544592 59027
rect 544018 58907 544508 58943
rect 543934 58823 544424 58859
rect 543850 58739 544340 58775
rect 543766 58655 544256 58691
rect 543682 58571 544172 58607
rect 543598 58487 544088 58523
rect 543514 58403 544004 58439
rect 543430 58319 543920 58355
rect 543346 58235 543836 58271
rect 543262 58151 543752 58187
rect 543178 58067 543668 58103
rect 543094 57983 543584 58019
rect 543010 57899 543500 57935
rect 542926 57815 543416 57851
rect 542842 57731 543332 57767
rect 542758 57647 543248 57683
rect 542674 57563 543164 57599
rect 542590 57479 543080 57515
rect 542506 57395 542996 57431
rect 542422 57311 542912 57347
rect 542338 57227 542828 57263
rect 542254 57143 542744 57179
rect 542170 57059 542660 57095
rect 542086 56975 542576 57011
rect 542002 56891 542492 56927
rect 541918 56807 542408 56843
rect 541834 56723 542324 56759
rect 541750 56639 542240 56675
rect 541666 56555 542156 56591
rect 541582 56471 542072 56507
rect 541175 54764 541731 55736
rect 541177 51312 541733 52284
rect 542036 50644 542072 56471
rect 540951 50608 542072 50644
rect 540268 49920 540338 49930
rect 540164 49836 540216 49842
rect 540164 49778 540216 49784
rect 540052 49751 540104 49757
rect 540052 49693 540104 49699
rect 534785 47953 535757 47959
rect 534885 47671 535757 47953
rect 534785 46968 535757 47671
rect 538237 46909 539209 47448
rect 528646 45792 530302 45828
rect 528562 45708 530218 45744
rect 528478 45624 530134 45660
rect 528394 45540 530050 45576
rect 528310 45456 529966 45492
rect 528226 45372 529882 45408
rect 528142 45288 529798 45324
rect 528058 45204 529714 45240
rect 527974 45120 529630 45156
rect 527890 45036 529546 45072
rect 527806 44952 529462 44988
rect 527722 44868 529378 44904
rect 527422 43866 529086 43902
rect 527350 43794 529000 43830
rect 527278 43722 528916 43758
rect 527206 43650 528832 43686
rect 527134 43578 528748 43614
rect 527062 43506 528664 43542
rect 526990 43434 528580 43470
rect 526918 43362 528496 43398
rect 526846 43290 528412 43326
rect 526774 43218 528328 43254
rect 526702 43146 528244 43182
rect 526630 43074 528160 43110
rect 526558 43002 528076 43038
rect 526486 42930 527992 42966
rect 526414 42858 527908 42894
rect 526342 42786 527824 42822
rect 526270 42714 527740 42750
rect 526198 42642 527656 42678
rect 526126 42570 527573 42606
rect 526054 42498 527488 42534
rect 525982 42426 527405 42462
rect 525910 42354 527320 42390
rect 525838 42282 527236 42318
rect 525766 42210 527153 42246
rect 525694 42138 527068 42174
rect 525622 42066 526984 42102
rect 525550 41994 526900 42030
rect 525478 41922 526816 41958
rect 525406 41850 526732 41886
rect 525334 41778 526648 41814
rect 525262 41706 526564 41742
rect 525190 41634 526480 41670
rect 525118 41562 526396 41598
rect 525046 41490 526312 41526
rect 524974 41418 526228 41454
rect 524902 41346 526146 41382
rect 524830 41274 526062 41310
rect 524758 41202 525978 41238
rect 524686 41130 525894 41166
rect 524614 41058 525810 41094
rect 524542 40986 525726 41022
rect 524470 40914 525642 40950
rect 524398 40842 525558 40878
rect 524326 40770 525474 40806
rect 524254 40698 525390 40734
rect 524182 40626 525306 40662
rect 524110 40554 525222 40590
rect 524038 40482 525138 40518
rect 523966 40410 525054 40446
rect 523894 40338 524970 40374
rect 523822 40266 524886 40302
rect 523750 40194 524802 40230
rect 523678 40122 524718 40158
rect 523510 37474 524462 37510
rect 523426 37390 524378 37426
rect 523342 37306 524294 37342
rect 523258 37222 524210 37258
rect 523174 37138 524126 37174
rect 523090 37054 524042 37090
rect 523006 36970 523958 37006
rect 522922 36886 523874 36922
rect 522838 36802 523790 36838
rect 522754 36718 523706 36754
rect 522670 36634 523622 36670
rect 522586 36550 523538 36586
rect 522502 36466 523454 36502
rect 522418 36382 523370 36418
rect 522035 27103 522999 27139
rect 521951 27019 522915 27055
rect 521867 26935 522831 26971
rect 521783 26851 522747 26887
rect 521699 26767 522663 26803
rect 521615 26683 522579 26719
rect 521530 26599 522495 26635
rect 521446 26515 522411 26551
rect 521362 26431 522327 26467
rect 521278 26347 522243 26383
rect 521194 26263 522159 26299
rect 521110 26179 522075 26215
rect 521026 26095 521991 26131
rect 520942 26011 521907 26047
rect 520858 25927 521823 25963
rect 520774 25843 521739 25879
rect 431742 22602 439077 22807
rect 431742 21785 431923 22602
rect 438850 21785 439077 22602
rect 472975 22662 478554 22814
rect 431742 21603 439077 21785
rect 464419 21999 464585 22012
rect 464419 21538 464430 21999
rect 464574 21538 464585 21999
rect 464419 21526 464585 21538
rect 464711 21998 464877 22012
rect 464711 21537 464722 21998
rect 464866 21537 464877 21998
rect 464711 21526 464877 21537
rect 465015 21997 465181 22012
rect 465015 21536 465027 21997
rect 465171 21536 465181 21997
rect 465015 21526 465181 21536
rect 465352 22001 465518 22013
rect 465352 21540 465360 22001
rect 465504 21540 465518 22001
rect 465352 21527 465518 21540
rect 467417 22000 467624 22011
rect 467417 21539 467428 22000
rect 467613 21539 467624 22000
rect 464477 20967 464513 21526
rect 464778 21053 464814 21526
rect 465074 21134 465110 21526
rect 465406 21219 465442 21527
rect 467417 21526 467624 21539
rect 472975 21637 473177 22662
rect 478353 21637 478554 22662
rect 467488 21305 467524 21526
rect 472975 21503 478554 21637
rect 467480 21299 467532 21305
rect 467480 21241 467532 21247
rect 465398 21213 465450 21219
rect 465398 21155 465450 21161
rect 465066 21128 465118 21134
rect 465066 21070 465118 21076
rect 464770 21047 464822 21053
rect 464770 20989 464822 20995
rect 464469 20961 464521 20967
rect 464469 20903 464521 20909
rect 482504 20002 482540 20018
rect 482496 19996 482548 20002
rect 482496 19938 482548 19944
rect 482420 19918 482456 19930
rect 482412 19912 482464 19918
rect 482412 19854 482464 19860
rect 482336 19834 482372 19846
rect 482328 19828 482380 19834
rect 482328 19770 482380 19776
rect 482252 19750 482288 19762
rect 482244 19744 482296 19750
rect 367620 19696 367737 19701
rect 367616 19589 367625 19696
rect 367732 19589 367741 19696
rect 482244 19686 482296 19692
rect 482168 19666 482204 19678
rect 482160 19660 482212 19666
rect 482160 19602 482212 19608
rect 354364 19356 354416 19362
rect 354364 19298 354416 19304
rect 354280 19272 354332 19278
rect 354280 19214 354332 19220
rect 354196 19188 354248 19194
rect 354196 19130 354248 19136
rect 354112 19104 354164 19110
rect 354112 19046 354164 19052
rect 354028 19020 354080 19026
rect 354028 18962 354080 18968
rect 353944 18936 353996 18942
rect 353944 18878 353996 18884
rect 353860 18852 353912 18858
rect 353860 18794 353912 18800
rect 353776 18768 353828 18774
rect 353776 18710 353828 18716
rect 353692 18684 353744 18690
rect 353692 18626 353744 18632
rect 353608 18600 353660 18606
rect 353608 18542 353660 18548
rect 353524 18516 353576 18522
rect 353524 18458 353576 18464
rect 353392 18432 353444 18438
rect 353392 18374 353444 18380
rect 353272 18264 353324 18270
rect 353272 18206 353324 18212
rect 353188 18180 353240 18186
rect 353188 18122 353240 18128
rect 353104 18096 353156 18102
rect 353104 18038 353156 18044
rect 353020 18012 353072 18018
rect 353020 17954 353072 17960
rect 352936 17928 352988 17934
rect 352936 17870 352988 17876
rect 352852 17844 352904 17850
rect 352852 17786 352904 17792
rect 352768 17760 352820 17766
rect 352768 17702 352820 17708
rect 352684 17676 352736 17682
rect 352684 17618 352736 17624
rect 353400 17510 353436 18374
rect 353392 17504 353444 17510
rect 353392 17446 353444 17452
rect 294461 16310 295062 16433
rect 367620 16297 367737 19589
rect 482084 19582 482120 19594
rect 482076 19576 482128 19582
rect 482076 19518 482128 19524
rect 482000 19498 482036 19510
rect 481992 19492 482044 19498
rect 481992 19434 482044 19440
rect 481916 19414 481952 19426
rect 481908 19408 481960 19414
rect 481908 19350 481960 19356
rect 481832 19330 481868 19342
rect 481824 19324 481876 19330
rect 481824 19266 481876 19272
rect 481748 19246 481784 19258
rect 481740 19240 481792 19246
rect 481740 19182 481792 19188
rect 481664 19162 481700 19174
rect 481656 19156 481708 19162
rect 481656 19098 481708 19104
rect 481580 19078 481616 19090
rect 481572 19072 481624 19078
rect 481572 19014 481624 19020
rect 481496 18994 481532 19006
rect 481488 18988 481540 18994
rect 481488 18930 481540 18936
rect 481412 18910 481448 18922
rect 481404 18904 481456 18910
rect 481404 18846 481456 18852
rect 481328 18826 481364 18838
rect 481320 18820 481372 18826
rect 481320 18762 481372 18768
rect 481244 18742 481280 18754
rect 481236 18736 481288 18742
rect 481236 18678 481288 18684
rect 481160 18658 481196 18670
rect 481152 18652 481204 18658
rect 481152 18594 481204 18600
rect 481076 18574 481112 18586
rect 481068 18568 481120 18574
rect 481068 18510 481120 18516
rect 480992 18490 481028 18502
rect 480984 18484 481036 18490
rect 480984 18426 481036 18432
rect 480908 18406 480944 18418
rect 480900 18400 480952 18406
rect 480900 18342 480952 18348
rect 480824 18322 480860 18334
rect 480816 18316 480868 18322
rect 480816 18258 480868 18264
rect 367620 16180 368062 16297
rect 367945 15849 368062 16180
rect 367945 15726 368062 15732
rect 480824 15286 480860 18258
rect 480908 15370 480944 18342
rect 480992 15454 481028 18426
rect 481076 15538 481112 18510
rect 481160 15622 481196 18594
rect 481244 15706 481280 18678
rect 481328 15790 481364 18762
rect 481412 15874 481448 18846
rect 481496 15958 481532 18930
rect 481580 16042 481616 19014
rect 481664 16126 481700 19098
rect 481748 16210 481784 19182
rect 481832 16294 481868 19266
rect 481916 16378 481952 19350
rect 482000 16462 482036 19434
rect 482084 16546 482120 19518
rect 482168 16630 482204 19602
rect 482252 16714 482288 19686
rect 482336 16798 482372 19770
rect 482420 16882 482456 19854
rect 482504 16966 482540 19938
rect 482504 16930 484736 16966
rect 482420 16846 484652 16882
rect 482336 16762 484568 16798
rect 482252 16678 484484 16714
rect 482168 16594 484400 16630
rect 482084 16510 484316 16546
rect 482000 16426 484232 16462
rect 481916 16342 484148 16378
rect 481832 16258 484064 16294
rect 481748 16174 483980 16210
rect 481664 16090 483896 16126
rect 481580 16006 483812 16042
rect 481496 15922 483728 15958
rect 481412 15838 483644 15874
rect 481328 15754 483560 15790
rect 481244 15670 483476 15706
rect 481160 15586 483392 15622
rect 481076 15502 483308 15538
rect 480992 15418 483224 15454
rect 480908 15334 483140 15370
rect 480824 15250 483056 15286
rect 363194 13545 363246 13551
rect 363194 13487 363246 13493
rect 290025 5332 290077 5338
rect 290025 5274 290077 5280
rect 289941 5248 289993 5254
rect 289941 5190 289993 5196
rect 289857 5164 289909 5170
rect 289857 5106 289909 5112
rect 289773 5080 289825 5086
rect 289773 5022 289825 5028
rect 289689 4996 289741 5002
rect 289689 4938 289741 4944
rect 289605 4912 289657 4918
rect 289605 4854 289657 4860
rect 289521 4828 289573 4834
rect 289521 4770 289573 4776
rect 289437 4744 289489 4750
rect 289437 4686 289489 4692
rect 289353 4660 289405 4666
rect 289353 4602 289405 4608
rect 289269 4576 289321 4582
rect 289269 4518 289321 4524
rect 289185 4492 289237 4498
rect 289185 4434 289237 4440
rect 289101 4408 289153 4414
rect 289101 4350 289153 4356
rect 289017 4324 289069 4330
rect 289017 4266 289069 4272
rect 288933 4240 288985 4246
rect 288933 4182 288985 4188
rect 288849 4156 288901 4162
rect 288849 4098 288901 4104
rect 288765 4072 288817 4078
rect 288765 4014 288817 4020
rect 288681 3988 288733 3994
rect 288681 3930 288733 3936
rect 288597 3904 288649 3910
rect 288597 3846 288649 3852
rect 288513 3820 288565 3826
rect 288513 3762 288565 3768
rect 288429 3736 288481 3742
rect 288429 3678 288481 3684
rect 288345 3652 288397 3658
rect 288345 3594 288397 3600
rect 288261 3568 288313 3574
rect 288261 3510 288313 3516
rect 288177 3484 288229 3490
rect 288177 3426 288229 3432
rect 288093 3400 288145 3406
rect 288093 3342 288145 3348
rect 288009 3316 288061 3322
rect 288009 3258 288061 3264
rect 287925 3232 287977 3238
rect 287925 3174 287977 3180
rect 287841 3148 287893 3154
rect 287841 3090 287893 3096
rect 287757 3064 287809 3070
rect 287757 3006 287809 3012
rect 287765 3000 287801 3006
rect 363201 2940 363237 13487
rect 363285 11921 363321 11930
rect 363280 11915 363332 11921
rect 363280 11857 363332 11863
rect 363196 2934 363248 2940
rect 363196 2876 363248 2882
rect 363201 2866 363237 2876
rect 286641 2375 286693 2381
rect 286641 2317 286693 2323
rect 273652 1426 273704 1432
rect 273652 1368 273704 1374
rect 273660 1367 273696 1368
rect 363285 504 363321 11857
rect 466898 2604 466938 7626
rect 467022 2688 467062 7626
rect 467138 2772 467178 7626
rect 467258 2856 467298 7626
rect 467249 2850 467301 2856
rect 467249 2792 467301 2798
rect 467258 2788 467298 2792
rect 467128 2766 467180 2772
rect 467128 2708 467180 2714
rect 467138 2703 467178 2708
rect 467015 2682 467067 2688
rect 467015 2624 467067 2630
rect 467022 2619 467062 2624
rect 466894 2598 466946 2604
rect 466894 2540 466946 2546
rect 466898 2535 466938 2540
rect 469490 2352 469530 7626
rect 469610 2436 469650 7626
rect 469603 2430 469655 2436
rect 469603 2372 469655 2378
rect 469610 2367 469650 2372
rect 469480 2346 469532 2352
rect 469480 2288 469532 2294
rect 469490 2285 469530 2288
rect 469730 1512 469770 7626
rect 469850 2520 469890 7626
rect 469841 2514 469893 2520
rect 469841 2456 469893 2462
rect 469850 2452 469890 2456
rect 472082 2016 472122 7626
rect 472202 2100 472242 7626
rect 472322 2268 472362 7626
rect 472313 2262 472365 2268
rect 472313 2202 472365 2210
rect 472442 2184 472482 7626
rect 472437 2178 472489 2184
rect 472437 2120 472489 2126
rect 472191 2094 472243 2100
rect 472191 2036 472243 2042
rect 472202 2034 472242 2036
rect 472073 2010 472125 2016
rect 472073 1952 472125 1958
rect 472082 1947 472122 1952
rect 474674 1680 474714 7626
rect 474794 1764 474834 7626
rect 474914 1932 474954 7626
rect 474907 1926 474959 1932
rect 474907 1868 474959 1874
rect 475034 1848 475074 7626
rect 475028 1842 475080 1848
rect 475028 1784 475080 1790
rect 475034 1778 475074 1784
rect 474785 1758 474837 1764
rect 474785 1700 474837 1706
rect 474794 1695 474834 1700
rect 474664 1674 474716 1680
rect 474664 1616 474716 1622
rect 474674 1611 474714 1616
rect 469722 1506 469774 1512
rect 469722 1448 469774 1454
rect 469730 1445 469770 1448
rect 477266 1092 477306 7626
rect 477386 1176 477426 7626
rect 477506 1596 477546 7626
rect 477498 1590 477550 1596
rect 477498 1532 477550 1538
rect 477506 1522 477546 1532
rect 477626 1260 477666 7626
rect 477614 1254 477666 1260
rect 477614 1196 477666 1202
rect 477626 1188 477666 1196
rect 477379 1170 477431 1176
rect 477379 1112 477431 1118
rect 477386 1105 477426 1112
rect 477258 1086 477310 1092
rect 477258 1028 477310 1034
rect 477266 1011 477306 1028
rect 479858 588 479898 7626
rect 479978 672 480018 7626
rect 480098 840 480138 7626
rect 480091 834 480143 840
rect 480091 776 480143 782
rect 480098 773 480138 776
rect 480218 756 480258 7626
rect 482450 1008 482490 7626
rect 482570 1344 482610 7626
rect 482561 1338 482613 1344
rect 482561 1280 482613 1286
rect 482570 1275 482610 1280
rect 482445 1002 482497 1008
rect 482445 944 482497 950
rect 482450 935 482490 944
rect 482690 924 482730 7626
rect 482810 1422 482850 7626
rect 483020 6858 483056 15250
rect 483104 6942 483140 15334
rect 483188 7026 483224 15418
rect 483272 7110 483308 15502
rect 483356 7194 483392 15586
rect 483440 7278 483476 15670
rect 483524 7362 483560 15754
rect 483608 7446 483644 15838
rect 483692 7530 483728 15922
rect 483776 7614 483812 16006
rect 483860 7698 483896 16090
rect 483944 7782 483980 16174
rect 484028 7866 484064 16258
rect 484112 7950 484148 16342
rect 484196 8034 484232 16426
rect 484280 8118 484316 16510
rect 484364 8202 484400 16594
rect 484448 8286 484484 16678
rect 484532 8370 484568 16762
rect 484616 8454 484652 16846
rect 484700 8538 484736 16930
rect 521026 14222 521032 14228
rect 520484 14182 521032 14222
rect 521026 14176 521032 14182
rect 521084 14176 521090 14228
rect 520942 14098 520948 14104
rect 520492 14058 520948 14098
rect 520942 14052 520948 14058
rect 521000 14052 521006 14104
rect 520854 13982 520860 13988
rect 520492 13942 520860 13982
rect 520854 13936 520860 13942
rect 520912 13936 520918 13988
rect 520770 13862 520776 13868
rect 520500 13822 520776 13862
rect 520770 13816 520776 13822
rect 520828 13816 520834 13868
rect 520692 11630 520698 11636
rect 490681 9730 490687 9798
rect 490755 9730 490761 9798
rect 484692 8532 484744 8538
rect 484692 8474 484744 8480
rect 484700 8470 484736 8474
rect 484608 8448 484660 8454
rect 484608 8390 484660 8396
rect 484616 8384 484652 8390
rect 484524 8364 484576 8370
rect 484524 8306 484576 8312
rect 484532 8304 484568 8306
rect 484440 8280 484492 8286
rect 484440 8222 484492 8228
rect 484448 8218 484484 8222
rect 484356 8196 484408 8202
rect 484356 8138 484408 8144
rect 484364 8132 484400 8138
rect 484272 8112 484324 8118
rect 484272 8054 484324 8060
rect 484280 8048 484316 8054
rect 484188 8028 484240 8034
rect 484188 7970 484240 7976
rect 484196 7964 484232 7970
rect 484104 7944 484156 7950
rect 484104 7886 484156 7892
rect 484112 7884 484148 7886
rect 484020 7860 484072 7866
rect 484020 7802 484072 7808
rect 484028 7796 484064 7802
rect 483936 7776 483988 7782
rect 483936 7718 483988 7724
rect 483944 7716 483980 7718
rect 483852 7692 483904 7698
rect 483852 7634 483904 7640
rect 483860 7632 483896 7634
rect 483768 7608 483820 7614
rect 483768 7550 483820 7556
rect 483684 7524 483736 7530
rect 483684 7466 483736 7472
rect 483692 7462 483728 7466
rect 483600 7440 483652 7446
rect 483600 7382 483652 7388
rect 483608 7378 483644 7382
rect 483516 7356 483568 7362
rect 483516 7298 483568 7304
rect 483524 7296 483560 7298
rect 483432 7272 483484 7278
rect 483432 7214 483484 7220
rect 483348 7188 483400 7194
rect 483348 7130 483400 7136
rect 483356 7128 483392 7130
rect 483264 7104 483316 7110
rect 483264 7046 483316 7052
rect 483272 7044 483308 7046
rect 483180 7020 483232 7026
rect 483180 6960 483232 6968
rect 483096 6936 483148 6942
rect 483096 6878 483148 6884
rect 483012 6852 483064 6858
rect 483012 6794 483064 6800
rect 490687 2938 490755 9730
rect 492916 7712 493066 11624
rect 520506 11590 520698 11630
rect 520692 11584 520698 11590
rect 520750 11584 520756 11636
rect 520606 11510 520612 11516
rect 520500 11470 520612 11510
rect 520606 11464 520612 11470
rect 520664 11464 520670 11516
rect 520520 11390 520526 11396
rect 520502 11350 520526 11390
rect 520520 11344 520526 11350
rect 520578 11344 520584 11396
rect 520436 11270 520442 11276
rect 520306 11230 520442 11270
rect 520436 11224 520442 11230
rect 520494 11224 520500 11276
rect 521703 8676 521739 25843
rect 521787 8760 521823 25927
rect 521871 8844 521907 26011
rect 521955 8928 521991 26095
rect 522039 9012 522075 26179
rect 522123 9096 522159 26263
rect 522207 9180 522243 26347
rect 522291 9264 522327 26431
rect 522375 9348 522411 26515
rect 522459 9432 522495 26599
rect 522543 9516 522579 26683
rect 522627 9600 522663 26767
rect 522711 9684 522747 26851
rect 522795 9768 522831 26935
rect 522879 9852 522915 27019
rect 522963 9936 522999 27103
rect 523334 14752 523370 36382
rect 523418 14836 523454 36466
rect 523502 14920 523538 36550
rect 523586 15004 523622 36634
rect 523670 15088 523706 36718
rect 523754 15172 523790 36802
rect 523838 15256 523874 36886
rect 523922 15340 523958 36970
rect 524006 15424 524042 37054
rect 524090 15508 524126 37138
rect 524174 15592 524210 37222
rect 524258 15676 524294 37306
rect 524342 15760 524378 37390
rect 524426 15844 524462 37474
rect 524418 15838 524470 15844
rect 524418 15780 524470 15786
rect 524334 15754 524386 15760
rect 524334 15696 524386 15702
rect 524250 15670 524302 15676
rect 524250 15612 524302 15618
rect 524166 15586 524218 15592
rect 524166 15528 524218 15534
rect 524082 15502 524134 15508
rect 524082 15444 524134 15450
rect 523998 15418 524050 15424
rect 523998 15360 524050 15366
rect 523914 15334 523966 15340
rect 523914 15276 523966 15282
rect 523830 15250 523882 15256
rect 523830 15192 523882 15198
rect 523746 15166 523798 15172
rect 523746 15108 523798 15114
rect 523662 15082 523714 15088
rect 523662 15024 523714 15030
rect 523578 14998 523630 15004
rect 523578 14940 523630 14946
rect 523494 14914 523546 14920
rect 523494 14856 523546 14862
rect 523410 14830 523462 14836
rect 523410 14772 523462 14778
rect 523326 14746 523378 14752
rect 523326 14688 523378 14694
rect 524682 10602 524718 40122
rect 524766 10676 524802 40194
rect 524850 10750 524886 40266
rect 524934 10824 524970 40338
rect 525018 10898 525054 40410
rect 525102 10972 525138 40482
rect 525186 11046 525222 40554
rect 525270 11120 525306 40626
rect 525354 11194 525390 40698
rect 525438 11268 525474 40770
rect 525522 11342 525558 40842
rect 525606 11416 525642 40914
rect 525690 11490 525726 40986
rect 525774 11564 525810 41058
rect 525858 11638 525894 41130
rect 525942 11712 525978 41202
rect 526026 11786 526062 41274
rect 526110 11860 526146 41346
rect 526192 11934 526228 41418
rect 526276 12008 526312 41490
rect 526360 12082 526396 41562
rect 526444 12156 526480 41634
rect 526528 12230 526564 41706
rect 526612 12304 526648 41778
rect 526696 12378 526732 41850
rect 526780 12452 526816 41922
rect 526864 12526 526900 41994
rect 526948 12600 526984 42066
rect 527032 12674 527068 42138
rect 527116 12748 527152 42210
rect 527200 12822 527236 42282
rect 527284 12896 527320 42354
rect 527368 12970 527404 42426
rect 527452 13044 527488 42498
rect 527536 13118 527572 42570
rect 527620 13192 527656 42642
rect 527704 13266 527740 42714
rect 527788 13340 527824 42786
rect 527872 13414 527908 42858
rect 527956 13488 527992 42930
rect 528040 13562 528076 43002
rect 528124 13636 528160 43074
rect 528208 13710 528244 43146
rect 528292 13784 528328 43218
rect 528376 13858 528412 43290
rect 528460 13932 528496 43362
rect 528544 14006 528580 43434
rect 528628 14080 528664 43506
rect 528712 14154 528748 43578
rect 528796 14228 528832 43650
rect 528880 14302 528916 43722
rect 528964 14376 529000 43794
rect 529048 39762 529086 43866
rect 529048 14450 529084 39762
rect 529342 17449 529378 44868
rect 529426 17533 529462 44952
rect 529510 17617 529546 45036
rect 529594 17701 529630 45120
rect 529678 17785 529714 45204
rect 529762 17869 529798 45288
rect 529846 17953 529882 45372
rect 529930 18037 529966 45456
rect 530014 18121 530050 45540
rect 530098 18205 530134 45624
rect 530182 18289 530218 45708
rect 530266 18373 530302 45792
rect 534785 34315 535755 34623
rect 538237 34221 539207 34639
rect 538208 33906 539207 34221
rect 538208 33426 539180 33906
rect 530464 21355 530492 21361
rect 530452 21349 530504 21355
rect 530452 21291 530504 21297
rect 530258 18367 530310 18373
rect 530258 18309 530310 18315
rect 530266 18304 530302 18309
rect 530174 18283 530226 18289
rect 530174 18225 530226 18231
rect 530182 18220 530218 18225
rect 530090 18199 530142 18205
rect 530090 18141 530142 18147
rect 530098 18136 530134 18141
rect 530006 18115 530058 18121
rect 530006 18057 530058 18063
rect 530014 18052 530050 18057
rect 529922 18031 529974 18037
rect 529922 17973 529974 17979
rect 529930 17968 529966 17973
rect 529838 17947 529890 17953
rect 529838 17889 529890 17895
rect 529846 17884 529882 17889
rect 529754 17863 529806 17869
rect 529754 17805 529806 17811
rect 529762 17800 529798 17805
rect 529670 17779 529722 17785
rect 529670 17721 529722 17727
rect 529678 17716 529714 17721
rect 529586 17695 529638 17701
rect 529586 17637 529638 17643
rect 529594 17632 529630 17637
rect 529502 17611 529554 17617
rect 529502 17553 529554 17559
rect 529510 17548 529546 17553
rect 529418 17527 529470 17533
rect 529418 17469 529470 17475
rect 529426 17464 529462 17469
rect 529334 17443 529386 17449
rect 529334 17385 529386 17391
rect 529342 17380 529378 17385
rect 529042 14444 529094 14450
rect 529042 14386 529094 14392
rect 529048 14382 529084 14386
rect 528958 14370 529010 14376
rect 528958 14312 529010 14318
rect 528964 14308 529000 14312
rect 528874 14296 528926 14302
rect 528874 14238 528926 14244
rect 528880 14234 528916 14238
rect 528790 14222 528842 14228
rect 528790 14164 528842 14170
rect 528796 14160 528832 14164
rect 528706 14148 528758 14154
rect 528706 14090 528758 14096
rect 528712 14086 528748 14090
rect 528622 14074 528674 14080
rect 528622 14016 528674 14022
rect 528628 14012 528664 14016
rect 528538 14000 528590 14006
rect 528538 13942 528590 13948
rect 528544 13938 528580 13942
rect 528454 13926 528506 13932
rect 528454 13868 528506 13874
rect 528460 13864 528496 13868
rect 528370 13852 528422 13858
rect 528370 13794 528422 13800
rect 528376 13790 528412 13794
rect 528286 13778 528338 13784
rect 528286 13720 528338 13726
rect 528292 13716 528328 13720
rect 528202 13704 528254 13710
rect 528202 13646 528254 13652
rect 528208 13642 528244 13646
rect 528118 13630 528170 13636
rect 528118 13572 528170 13578
rect 528124 13568 528160 13572
rect 528034 13556 528086 13562
rect 528034 13498 528086 13504
rect 528040 13494 528076 13498
rect 527950 13482 528002 13488
rect 527950 13424 528002 13430
rect 527956 13420 527992 13424
rect 527866 13408 527918 13414
rect 527866 13350 527918 13356
rect 527872 13346 527908 13350
rect 527782 13334 527834 13340
rect 527782 13276 527834 13282
rect 527788 13272 527824 13276
rect 527698 13260 527750 13266
rect 527698 13202 527750 13208
rect 527704 13198 527740 13202
rect 527614 13186 527666 13192
rect 527614 13128 527666 13134
rect 527620 13124 527656 13128
rect 527530 13112 527582 13118
rect 527530 13054 527582 13060
rect 527536 13050 527572 13054
rect 527446 13038 527498 13044
rect 527446 12980 527498 12986
rect 527452 12976 527488 12980
rect 527362 12964 527414 12970
rect 527362 12906 527414 12912
rect 527368 12902 527404 12906
rect 527278 12890 527330 12896
rect 527278 12832 527330 12838
rect 527284 12828 527320 12832
rect 527194 12816 527246 12822
rect 527194 12758 527246 12764
rect 527200 12754 527236 12758
rect 527110 12742 527162 12748
rect 527110 12684 527162 12690
rect 527116 12680 527152 12684
rect 527026 12668 527078 12674
rect 527026 12610 527078 12616
rect 527032 12606 527068 12610
rect 526942 12594 526994 12600
rect 526942 12536 526994 12542
rect 526948 12532 526984 12536
rect 526858 12520 526910 12526
rect 526858 12462 526910 12468
rect 526864 12458 526900 12462
rect 526774 12446 526826 12452
rect 526774 12388 526826 12394
rect 526780 12384 526816 12388
rect 526690 12372 526742 12378
rect 526690 12314 526742 12320
rect 526696 12310 526732 12314
rect 526606 12298 526658 12304
rect 526606 12240 526658 12246
rect 526612 12236 526648 12240
rect 526522 12224 526574 12230
rect 526522 12166 526574 12172
rect 526528 12162 526564 12166
rect 526438 12150 526490 12156
rect 526438 12092 526490 12098
rect 526444 12088 526480 12092
rect 526354 12076 526406 12082
rect 526354 12018 526406 12024
rect 530464 12020 530492 21291
rect 530548 21271 530576 21277
rect 530536 21265 530588 21271
rect 530536 21207 530588 21213
rect 526360 12014 526396 12018
rect 526270 12002 526322 12008
rect 526270 11944 526322 11950
rect 527520 11992 530492 12020
rect 526276 11940 526312 11944
rect 526186 11928 526238 11934
rect 526186 11870 526238 11876
rect 526192 11866 526228 11870
rect 526102 11854 526154 11860
rect 526102 11796 526154 11802
rect 526110 11792 526146 11796
rect 526018 11780 526070 11786
rect 526018 11722 526070 11728
rect 526026 11718 526062 11722
rect 525934 11706 525986 11712
rect 525934 11648 525986 11654
rect 525942 11644 525978 11648
rect 525850 11632 525902 11638
rect 525850 11574 525902 11580
rect 525858 11570 525894 11574
rect 525766 11558 525818 11564
rect 525766 11500 525818 11506
rect 525774 11496 525810 11500
rect 525682 11484 525734 11490
rect 525682 11426 525734 11432
rect 525690 11422 525726 11426
rect 525598 11410 525650 11416
rect 525598 11352 525650 11358
rect 525606 11348 525642 11352
rect 525514 11336 525566 11342
rect 525514 11278 525566 11284
rect 525522 11274 525558 11278
rect 525430 11262 525482 11268
rect 525430 11204 525482 11210
rect 525438 11200 525474 11204
rect 525346 11188 525398 11194
rect 525346 11130 525398 11136
rect 525354 11126 525390 11130
rect 525262 11114 525314 11120
rect 525262 11056 525314 11062
rect 525270 11052 525306 11056
rect 525178 11040 525230 11046
rect 525178 10982 525230 10988
rect 525186 10978 525222 10982
rect 525094 10966 525146 10972
rect 525094 10908 525146 10914
rect 525102 10904 525138 10908
rect 525010 10892 525062 10898
rect 525010 10834 525062 10840
rect 525018 10830 525054 10834
rect 524926 10818 524978 10824
rect 524926 10760 524978 10766
rect 524934 10756 524970 10760
rect 524842 10744 524894 10750
rect 524842 10686 524894 10692
rect 524850 10682 524886 10686
rect 524758 10670 524810 10676
rect 524758 10612 524810 10618
rect 524766 10608 524802 10612
rect 524674 10596 524726 10602
rect 524674 10538 524726 10544
rect 524682 10534 524718 10538
rect 522955 9930 523007 9936
rect 522955 9872 523007 9878
rect 522963 9870 522999 9872
rect 522871 9846 522923 9852
rect 522871 9788 522923 9794
rect 522879 9786 522915 9788
rect 522787 9762 522839 9768
rect 522787 9704 522839 9710
rect 522795 9702 522831 9704
rect 522703 9678 522755 9684
rect 522703 9620 522755 9626
rect 522711 9618 522747 9620
rect 522619 9594 522671 9600
rect 522619 9536 522671 9542
rect 522627 9534 522663 9536
rect 522535 9510 522587 9516
rect 522535 9452 522587 9458
rect 522543 9450 522579 9452
rect 522451 9426 522503 9432
rect 522451 9368 522503 9374
rect 522459 9366 522495 9368
rect 522367 9342 522419 9348
rect 522367 9284 522419 9290
rect 522375 9282 522411 9284
rect 522283 9258 522335 9264
rect 522283 9200 522335 9206
rect 522291 9198 522327 9200
rect 522199 9174 522251 9180
rect 522199 9116 522251 9122
rect 522207 9114 522243 9116
rect 522115 9090 522167 9096
rect 522115 9032 522167 9038
rect 522123 9030 522159 9032
rect 522031 9006 522083 9012
rect 522031 8948 522083 8954
rect 522039 8946 522075 8948
rect 521947 8922 521999 8928
rect 521947 8864 521999 8870
rect 521955 8862 521991 8864
rect 521863 8838 521915 8844
rect 521863 8780 521915 8786
rect 521871 8778 521907 8780
rect 521779 8754 521831 8760
rect 521779 8696 521831 8702
rect 521787 8694 521823 8696
rect 521695 8670 521747 8676
rect 521695 8612 521747 8618
rect 521703 8610 521739 8612
rect 490687 2864 490755 2870
rect 482798 1370 482804 1422
rect 482856 1370 482862 1422
rect 482810 1363 482850 1370
rect 482685 918 482737 924
rect 482685 860 482737 866
rect 482690 852 482730 860
rect 480207 750 480259 756
rect 480207 692 480259 698
rect 479966 666 480018 672
rect 479966 608 480018 614
rect 479978 599 480018 608
rect 479847 582 479899 588
rect 479847 524 479899 530
rect 479858 519 479898 524
rect 363277 498 363329 504
rect 363277 440 363329 446
rect 527520 0 527548 11992
rect 530548 11908 530576 21207
rect 530632 21187 530660 21193
rect 530620 21181 530672 21187
rect 530620 21123 530672 21129
rect 527632 11880 530576 11908
rect 527632 0 527660 11880
rect 530632 11796 530660 21123
rect 530716 21103 530744 21109
rect 530704 21097 530756 21103
rect 530704 21039 530756 21045
rect 527744 11768 530660 11796
rect 527744 0 527772 11768
rect 530716 11684 530744 21039
rect 530800 21019 530828 21025
rect 530788 21013 530840 21019
rect 530788 20955 530840 20961
rect 527856 11656 530744 11684
rect 527856 0 527884 11656
rect 530800 11572 530828 20955
rect 530884 20935 530912 20941
rect 530872 20929 530924 20935
rect 530872 20871 530924 20877
rect 527968 11544 530828 11572
rect 527968 0 527996 11544
rect 530884 11460 530912 20871
rect 530968 20851 530996 20857
rect 530956 20845 531008 20851
rect 530956 20787 531008 20793
rect 528080 11432 530912 11460
rect 528080 0 528108 11432
rect 530968 11348 530996 20787
rect 531052 20767 531080 20773
rect 531040 20761 531092 20767
rect 531040 20703 531092 20709
rect 528192 11320 530996 11348
rect 528192 0 528220 11320
rect 531052 11236 531080 20703
rect 531136 20683 531164 20689
rect 531124 20677 531176 20683
rect 531124 20619 531176 20625
rect 528304 11208 531080 11236
rect 528304 0 528332 11208
rect 531136 11124 531164 20619
rect 531220 20599 531248 20605
rect 531208 20593 531260 20599
rect 531208 20535 531260 20541
rect 528416 11096 531164 11124
rect 528416 0 528444 11096
rect 531220 11012 531248 20535
rect 534756 20522 535726 21104
rect 531304 20515 531332 20521
rect 531292 20509 531344 20515
rect 531292 20451 531344 20457
rect 528528 10984 531248 11012
rect 528528 0 528556 10984
rect 531304 10900 531332 20451
rect 531388 20431 531416 20437
rect 531376 20425 531428 20431
rect 531376 20367 531428 20373
rect 528640 10872 531332 10900
rect 528640 0 528668 10872
rect 531388 10788 531416 20367
rect 531472 20347 531500 20353
rect 531460 20341 531512 20347
rect 531460 20283 531512 20289
rect 528752 10760 531416 10788
rect 528752 0 528780 10760
rect 531472 10676 531500 20283
rect 531556 20263 531584 20269
rect 531544 20257 531596 20263
rect 531544 20199 531596 20205
rect 528864 10648 531500 10676
rect 528864 0 528892 10648
rect 531556 10564 531584 20199
rect 531640 20179 531668 20185
rect 531628 20173 531680 20179
rect 531628 20115 531680 20121
rect 538208 20150 539178 21257
rect 528976 10536 531584 10564
rect 528976 0 529004 10536
rect 531640 10452 531668 20115
rect 531724 20095 531752 20101
rect 531712 20089 531764 20095
rect 531712 20031 531764 20037
rect 529088 10424 531668 10452
rect 529088 0 529116 10424
rect 531724 10340 531752 20031
rect 531808 20011 531836 20017
rect 531796 20005 531848 20011
rect 531796 19947 531848 19953
rect 529200 10312 531752 10340
rect 529200 0 529228 10312
rect 531808 10228 531836 19947
rect 531892 19927 531920 19933
rect 531880 19921 531932 19927
rect 531880 19863 531932 19869
rect 529312 10200 531836 10228
rect 529312 0 529340 10200
rect 531892 10116 531920 19863
rect 531976 19843 532004 19849
rect 531964 19837 532016 19843
rect 531964 19779 532016 19785
rect 529424 10088 531920 10116
rect 529424 0 529452 10088
rect 531976 10004 532004 19779
rect 532060 19759 532088 19765
rect 532048 19753 532100 19759
rect 532048 19695 532100 19701
rect 529536 9976 532004 10004
rect 529536 0 529564 9976
rect 532060 9892 532088 19695
rect 532144 19675 532172 19681
rect 532132 19669 532184 19675
rect 532132 19611 532184 19617
rect 529648 9864 532088 9892
rect 529648 0 529676 9864
rect 532144 9780 532172 19611
rect 532228 19591 532256 19597
rect 532216 19585 532268 19591
rect 532216 19527 532268 19533
rect 529760 9752 532172 9780
rect 529760 0 529788 9752
rect 532228 9668 532256 19527
rect 532312 19507 532340 19513
rect 532300 19501 532352 19507
rect 532300 19443 532352 19449
rect 529872 9640 532256 9668
rect 529872 0 529900 9640
rect 532312 9556 532340 19443
rect 532396 19423 532424 19429
rect 532384 19417 532436 19423
rect 532384 19359 532436 19365
rect 529984 9528 532340 9556
rect 529984 0 530012 9528
rect 532396 9444 532424 19359
rect 532480 19339 532508 19345
rect 532468 19333 532520 19339
rect 532468 19275 532520 19281
rect 530096 9416 532424 9444
rect 530096 0 530124 9416
rect 532480 9332 532508 19275
rect 532564 19255 532592 19261
rect 532552 19249 532604 19255
rect 532552 19191 532604 19197
rect 530208 9304 532508 9332
rect 530208 0 530236 9304
rect 532564 9220 532592 19191
rect 538208 19181 539378 20150
rect 532648 19171 532676 19177
rect 532636 19165 532688 19171
rect 532636 19107 532688 19113
rect 530320 9192 532592 9220
rect 530320 0 530348 9192
rect 532648 9108 532676 19107
rect 532732 19087 532760 19093
rect 532720 19081 532772 19087
rect 532720 19023 532772 19029
rect 530432 9080 532676 9108
rect 530432 0 530460 9080
rect 532732 8996 532760 19023
rect 532816 19003 532844 19009
rect 532804 18997 532856 19003
rect 532804 18939 532856 18945
rect 530544 8968 532760 8996
rect 530544 0 530572 8968
rect 532816 8884 532844 18939
rect 532900 18919 532928 18925
rect 532888 18913 532940 18919
rect 532888 18855 532940 18861
rect 530656 8856 532844 8884
rect 530656 0 530684 8856
rect 532900 8772 532928 18855
rect 532984 18835 533012 18841
rect 532972 18829 533024 18835
rect 532972 18771 533024 18777
rect 530768 8744 532928 8772
rect 530768 0 530796 8744
rect 532984 8660 533012 18771
rect 533068 18751 533096 18757
rect 533056 18745 533108 18751
rect 533056 18687 533108 18693
rect 530880 8632 533012 8660
rect 530880 0 530908 8632
rect 533068 8548 533096 18687
rect 533152 18667 533180 18673
rect 533140 18661 533192 18667
rect 533140 18603 533192 18609
rect 530992 8520 533096 8548
rect 530992 0 531020 8520
rect 533152 8436 533180 18603
rect 533236 18583 533264 18589
rect 533224 18577 533276 18583
rect 533224 18519 533276 18525
rect 531104 8408 533180 8436
rect 531104 0 531132 8408
rect 533236 8324 533264 18519
rect 533320 18499 533348 18505
rect 533308 18493 533360 18499
rect 533308 18435 533360 18441
rect 531216 8296 533264 8324
rect 531216 0 531244 8296
rect 533320 8212 533348 18435
rect 538160 18372 538188 18375
rect 538148 18366 538200 18372
rect 538148 18308 538200 18314
rect 538048 18288 538076 18291
rect 538036 18282 538088 18288
rect 538036 18224 538088 18230
rect 537936 18204 537964 18207
rect 537924 18198 537976 18204
rect 537924 18140 537976 18146
rect 537824 18120 537852 18123
rect 537812 18114 537864 18120
rect 537812 18056 537864 18062
rect 537712 18036 537740 18039
rect 537700 18030 537752 18036
rect 537700 17972 537752 17978
rect 537600 17952 537628 17955
rect 537588 17946 537640 17952
rect 537588 17888 537640 17894
rect 537488 17868 537516 17871
rect 537476 17862 537528 17868
rect 537476 17804 537528 17810
rect 537376 17784 537404 17787
rect 537364 17778 537416 17784
rect 537364 17720 537416 17726
rect 537264 17700 537292 17703
rect 537252 17694 537304 17700
rect 537252 17636 537304 17642
rect 537152 17616 537180 17619
rect 537140 17610 537192 17616
rect 537140 17552 537192 17558
rect 537040 17532 537068 17535
rect 537028 17526 537080 17532
rect 537028 17468 537080 17474
rect 536928 17448 536956 17451
rect 536916 17442 536968 17448
rect 536916 17384 536968 17390
rect 536704 17138 536732 17148
rect 536692 17132 536744 17138
rect 536692 17074 536744 17080
rect 536592 17054 536620 17064
rect 536580 17048 536632 17054
rect 536580 16990 536632 16996
rect 536480 16970 536508 16980
rect 536468 16964 536520 16970
rect 536468 16906 536520 16912
rect 536368 16886 536396 16896
rect 536356 16880 536408 16886
rect 536356 16822 536408 16828
rect 536256 16802 536284 16812
rect 536244 16796 536296 16802
rect 536244 16738 536296 16744
rect 536144 16718 536172 16728
rect 536132 16712 536184 16718
rect 536132 16654 536184 16660
rect 536032 16634 536060 16644
rect 536020 16628 536072 16634
rect 536020 16570 536072 16576
rect 535920 16550 535948 16560
rect 535908 16544 535960 16550
rect 535908 16486 535960 16492
rect 535808 16466 535836 16476
rect 535796 16460 535848 16466
rect 535796 16402 535848 16408
rect 535696 16382 535724 16392
rect 535684 16376 535736 16382
rect 535684 16318 535736 16324
rect 535584 16298 535612 16308
rect 535572 16292 535624 16298
rect 535572 16234 535624 16240
rect 535472 16214 535500 16224
rect 535460 16208 535512 16214
rect 535460 16150 535512 16156
rect 535360 16130 535388 16140
rect 535348 16124 535400 16130
rect 535348 16066 535400 16072
rect 534800 10386 534828 10391
rect 534788 10380 534840 10386
rect 534788 10322 534840 10328
rect 531328 8184 533348 8212
rect 531328 0 531356 8184
rect 534688 2943 534716 2954
rect 534676 2937 534728 2943
rect 534676 2879 534728 2885
rect 534576 2859 534604 2870
rect 534564 2853 534616 2859
rect 534564 2795 534616 2801
rect 534464 2775 534492 2786
rect 534452 2769 534504 2775
rect 534452 2711 534504 2717
rect 534352 2691 534380 2702
rect 534340 2685 534392 2691
rect 534340 2627 534392 2633
rect 534240 2607 534268 2618
rect 534228 2601 534280 2607
rect 534228 2543 534280 2549
rect 534128 2523 534156 2534
rect 534116 2517 534168 2523
rect 534116 2459 534168 2465
rect 534016 2439 534044 2450
rect 534004 2433 534056 2439
rect 534004 2375 534056 2381
rect 533904 2355 533932 2366
rect 533892 2349 533944 2355
rect 533892 2291 533944 2297
rect 533792 2271 533820 2282
rect 533780 2265 533832 2271
rect 533780 2207 533832 2213
rect 533680 2187 533708 2198
rect 533668 2181 533720 2187
rect 533668 2123 533720 2129
rect 533568 2103 533596 2114
rect 533556 2097 533608 2103
rect 533556 2039 533608 2045
rect 533456 2019 533484 2030
rect 533444 2013 533496 2019
rect 533444 1955 533496 1961
rect 533344 1935 533372 1946
rect 533332 1929 533384 1935
rect 533332 1871 533384 1877
rect 533232 1851 533260 1862
rect 533220 1845 533272 1851
rect 533220 1787 533272 1793
rect 533120 1767 533148 1778
rect 533108 1761 533160 1767
rect 533108 1703 533160 1709
rect 533008 1683 533036 1694
rect 532996 1677 533048 1683
rect 532996 1619 533048 1625
rect 532896 1599 532924 1610
rect 532884 1593 532936 1599
rect 532884 1535 532936 1541
rect 532784 1515 532812 1526
rect 532772 1509 532824 1515
rect 532772 1451 532824 1457
rect 532672 1431 532700 1442
rect 532660 1425 532712 1431
rect 532660 1367 532712 1373
rect 532560 1347 532588 1358
rect 532548 1341 532600 1347
rect 532548 1283 532600 1289
rect 532448 1263 532476 1274
rect 532436 1257 532488 1263
rect 532436 1199 532488 1205
rect 532336 1179 532364 1190
rect 532324 1173 532376 1179
rect 532324 1115 532376 1121
rect 532224 1095 532252 1106
rect 532212 1089 532264 1095
rect 532212 1031 532264 1037
rect 532112 1011 532140 1022
rect 532100 1005 532152 1011
rect 532100 947 532152 953
rect 532000 927 532028 938
rect 531988 921 532040 927
rect 531988 863 532040 869
rect 531888 843 531916 854
rect 531876 837 531928 843
rect 531876 779 531928 785
rect 531776 759 531804 770
rect 531764 753 531816 759
rect 531764 695 531816 701
rect 531664 675 531692 686
rect 531652 669 531704 675
rect 531652 611 531704 617
rect 531552 591 531580 602
rect 531540 585 531592 591
rect 531540 527 531592 533
rect 531440 507 531468 518
rect 531428 501 531480 507
rect 531428 443 531480 449
rect 531440 0 531468 443
rect 531552 0 531580 527
rect 531664 0 531692 611
rect 531776 0 531804 695
rect 531888 0 531916 779
rect 532000 0 532028 863
rect 532112 0 532140 947
rect 532224 0 532252 1031
rect 532336 0 532364 1115
rect 532448 0 532476 1199
rect 532560 0 532588 1283
rect 532672 0 532700 1367
rect 532784 0 532812 1451
rect 532896 0 532924 1535
rect 533008 0 533036 1619
rect 533120 0 533148 1703
rect 533232 0 533260 1787
rect 533344 0 533372 1871
rect 533456 0 533484 1955
rect 533568 0 533596 2039
rect 533680 0 533708 2123
rect 533792 0 533820 2207
rect 533904 0 533932 2291
rect 534016 0 534044 2375
rect 534128 0 534156 2459
rect 534240 0 534268 2543
rect 534352 0 534380 2627
rect 534464 0 534492 2711
rect 534576 0 534604 2795
rect 534688 0 534716 2879
rect 534800 0 534828 10322
rect 535248 10295 535276 10310
rect 535230 10243 535236 10295
rect 535288 10243 535294 10295
rect 535136 10217 535164 10228
rect 535124 10211 535176 10217
rect 535124 10153 535176 10159
rect 535024 10133 535052 10141
rect 535012 10127 535064 10133
rect 535012 10069 535064 10075
rect 534912 10047 534940 10059
rect 534900 10041 534952 10047
rect 534900 9983 534952 9989
rect 534912 0 534940 9983
rect 535024 0 535052 10069
rect 535136 0 535164 10153
rect 535248 0 535276 10243
rect 535360 0 535388 16066
rect 535472 0 535500 16150
rect 535584 0 535612 16234
rect 535696 0 535724 16318
rect 535808 0 535836 16402
rect 535920 0 535948 16486
rect 536032 0 536060 16570
rect 536144 0 536172 16654
rect 536256 0 536284 16738
rect 536368 0 536396 16822
rect 536480 0 536508 16906
rect 536592 0 536620 16990
rect 536704 0 536732 17074
rect 536816 0 536844 350
rect 536928 0 536956 17384
rect 537040 0 537068 17468
rect 537152 0 537180 17552
rect 537264 0 537292 17636
rect 537376 0 537404 17720
rect 537488 0 537516 17804
rect 537600 0 537628 17888
rect 537712 0 537740 17972
rect 537824 0 537852 18056
rect 537936 0 537964 18140
rect 538048 0 538076 18224
rect 538160 0 538188 18308
rect 538408 16711 539378 19181
rect 539952 9938 539980 9948
rect 539940 9932 539992 9938
rect 539940 9874 539992 9880
rect 539840 9854 539868 9864
rect 539828 9848 539880 9854
rect 539828 9790 539880 9796
rect 539728 9770 539756 9780
rect 539716 9764 539768 9770
rect 539716 9706 539768 9712
rect 539616 9686 539644 9696
rect 539604 9680 539656 9686
rect 539604 9622 539656 9628
rect 539504 9602 539532 9612
rect 539492 9596 539544 9602
rect 539492 9538 539544 9544
rect 539392 9518 539420 9528
rect 539380 9512 539432 9518
rect 539380 9454 539432 9460
rect 539280 9434 539308 9444
rect 539268 9428 539320 9434
rect 539268 9370 539320 9376
rect 539168 9350 539196 9360
rect 539156 9344 539208 9350
rect 539156 9286 539208 9292
rect 539056 9266 539084 9276
rect 539044 9260 539096 9266
rect 539044 9202 539096 9208
rect 538944 9182 538972 9192
rect 538932 9176 538984 9182
rect 538932 9118 538984 9124
rect 538832 9098 538860 9108
rect 538820 9092 538872 9098
rect 538820 9034 538872 9040
rect 538720 9014 538748 9024
rect 538708 9008 538760 9014
rect 538708 8950 538760 8956
rect 538608 8930 538636 8940
rect 538596 8924 538648 8930
rect 538596 8866 538648 8872
rect 538496 8846 538524 8856
rect 538484 8840 538536 8846
rect 538484 8782 538536 8788
rect 538384 8762 538412 8772
rect 538372 8756 538424 8762
rect 538372 8698 538424 8704
rect 538272 8677 538300 8688
rect 538260 8671 538312 8677
rect 538260 8613 538312 8619
rect 538272 0 538300 8613
rect 538384 0 538412 8698
rect 538496 0 538524 8782
rect 538608 0 538636 8866
rect 538720 0 538748 8950
rect 538832 0 538860 9034
rect 538944 0 538972 9118
rect 539056 0 539084 9202
rect 539168 0 539196 9286
rect 539280 0 539308 9370
rect 539392 0 539420 9454
rect 539504 0 539532 9538
rect 539616 0 539644 9622
rect 539728 0 539756 9706
rect 539840 0 539868 9790
rect 539952 0 539980 9874
rect 540064 0 540092 49693
rect 540176 0 540204 49778
rect 540268 49693 540273 49920
rect 540332 49693 540338 49920
rect 540268 0 540338 49693
rect 540951 21355 540987 50608
rect 542120 50560 542156 56555
rect 541035 50524 542156 50560
rect 540943 21349 540995 21355
rect 540943 21291 540995 21297
rect 540951 21272 540987 21291
rect 541035 21271 541071 50524
rect 542204 50476 542240 56639
rect 541119 50440 542240 50476
rect 541027 21265 541079 21271
rect 541027 21207 541079 21213
rect 541035 21188 541071 21207
rect 541119 21187 541155 50440
rect 542288 50392 542324 56723
rect 541203 50356 542324 50392
rect 541111 21181 541163 21187
rect 541111 21123 541163 21129
rect 541119 21104 541155 21123
rect 541203 21103 541239 50356
rect 542372 50308 542408 56807
rect 541287 50272 542408 50308
rect 541195 21097 541247 21103
rect 541195 21039 541247 21045
rect 541203 21020 541239 21039
rect 541287 21019 541323 50272
rect 542456 50224 542492 56891
rect 541371 50188 542492 50224
rect 541279 21013 541331 21019
rect 541279 20955 541331 20961
rect 541287 20936 541323 20955
rect 541371 20935 541407 50188
rect 542540 50140 542576 56975
rect 541455 50104 542576 50140
rect 541363 20929 541415 20935
rect 541363 20871 541415 20877
rect 541371 20852 541407 20871
rect 541455 20851 541491 50104
rect 542624 50056 542660 57059
rect 541539 50020 542660 50056
rect 541447 20845 541499 20851
rect 541447 20787 541499 20793
rect 541455 20768 541491 20787
rect 541539 20767 541575 50020
rect 542708 49972 542744 57143
rect 541623 49936 542744 49972
rect 541531 20761 541583 20767
rect 541531 20703 541583 20709
rect 541539 20684 541575 20703
rect 541623 20683 541659 49936
rect 542792 49888 542828 57227
rect 541707 49852 542828 49888
rect 541615 20677 541667 20683
rect 541615 20619 541667 20625
rect 541623 20600 541659 20619
rect 541707 20599 541743 49852
rect 542876 49804 542912 57311
rect 541791 49768 542912 49804
rect 541699 20593 541751 20599
rect 541699 20535 541751 20541
rect 541707 20516 541743 20535
rect 541791 20515 541827 49768
rect 542960 49720 542996 57395
rect 541875 49684 542996 49720
rect 541783 20509 541835 20515
rect 541783 20451 541835 20457
rect 541791 20432 541827 20451
rect 541875 20431 541911 49684
rect 543044 49636 543080 57479
rect 541959 49600 543080 49636
rect 541867 20425 541919 20431
rect 541867 20367 541919 20373
rect 541875 20348 541911 20367
rect 541959 20347 541995 49600
rect 543128 49552 543164 57563
rect 542043 49516 543164 49552
rect 541951 20341 542003 20347
rect 541951 20283 542003 20289
rect 541959 20264 541995 20283
rect 542043 20263 542079 49516
rect 543212 49468 543248 57647
rect 542127 49432 543248 49468
rect 542035 20257 542087 20263
rect 542035 20199 542087 20205
rect 542043 20180 542079 20199
rect 542127 20179 542163 49432
rect 543296 49384 543332 57731
rect 542211 49348 543332 49384
rect 542119 20173 542171 20179
rect 542119 20115 542171 20121
rect 542127 20096 542163 20115
rect 542211 20095 542247 49348
rect 543380 49300 543416 57815
rect 542295 49264 543416 49300
rect 542203 20089 542255 20095
rect 542203 20031 542255 20037
rect 542211 20012 542247 20031
rect 542295 20011 542331 49264
rect 543464 49216 543500 57899
rect 542379 49180 543500 49216
rect 542287 20005 542339 20011
rect 542287 19947 542339 19953
rect 542295 19928 542331 19947
rect 542379 19927 542415 49180
rect 543548 49132 543584 57983
rect 542463 49096 543584 49132
rect 542371 19921 542423 19927
rect 542371 19863 542423 19869
rect 542379 19844 542415 19863
rect 542463 19843 542499 49096
rect 543632 49048 543668 58067
rect 542547 49012 543668 49048
rect 542455 19837 542507 19843
rect 542455 19779 542507 19785
rect 542463 19760 542499 19779
rect 542547 19759 542583 49012
rect 543716 48964 543752 58151
rect 542631 48928 543752 48964
rect 542539 19753 542591 19759
rect 542539 19695 542591 19701
rect 542547 19676 542583 19695
rect 542631 19675 542667 48928
rect 543800 48880 543836 58235
rect 542715 48844 543836 48880
rect 542623 19669 542675 19675
rect 542623 19611 542675 19617
rect 542631 19592 542667 19611
rect 542715 19591 542751 48844
rect 543884 48796 543920 58319
rect 542799 48760 543920 48796
rect 542707 19585 542759 19591
rect 542707 19527 542759 19533
rect 542715 19508 542751 19527
rect 542799 19507 542835 48760
rect 543968 48712 544004 58403
rect 542883 48676 544004 48712
rect 542791 19501 542843 19507
rect 542791 19443 542843 19449
rect 542799 19424 542835 19443
rect 542883 19423 542919 48676
rect 544052 48628 544088 58487
rect 542967 48592 544088 48628
rect 542875 19417 542927 19423
rect 542875 19359 542927 19365
rect 542883 19340 542919 19359
rect 542967 19339 543003 48592
rect 544136 48544 544172 58571
rect 543051 48508 544172 48544
rect 542959 19333 543011 19339
rect 542959 19275 543011 19281
rect 542967 19256 543003 19275
rect 543051 19255 543087 48508
rect 544220 48460 544256 58655
rect 543135 48424 544256 48460
rect 543043 19249 543095 19255
rect 543043 19191 543095 19197
rect 543051 19172 543087 19191
rect 543135 19171 543171 48424
rect 544304 48376 544340 58739
rect 543219 48340 544340 48376
rect 543127 19165 543179 19171
rect 543127 19107 543179 19113
rect 543135 19088 543171 19107
rect 543219 19087 543255 48340
rect 544388 48292 544424 58823
rect 543303 48256 544424 48292
rect 543211 19081 543263 19087
rect 543211 19023 543263 19029
rect 543219 19019 543255 19023
rect 543303 19003 543339 48256
rect 544472 48208 544508 58907
rect 543387 48172 544508 48208
rect 543295 18997 543347 19003
rect 543295 18939 543347 18945
rect 543303 18935 543339 18939
rect 543387 18919 543423 48172
rect 544556 48124 544592 58991
rect 543471 48088 544592 48124
rect 543379 18913 543431 18919
rect 543379 18855 543431 18861
rect 543387 18851 543423 18855
rect 543471 18835 543507 48088
rect 544640 48040 544676 59075
rect 543555 48004 544676 48040
rect 543463 18829 543515 18835
rect 543463 18771 543515 18777
rect 543471 18767 543507 18771
rect 543555 18751 543591 48004
rect 544724 47956 544760 59159
rect 543639 47920 544760 47956
rect 543547 18745 543599 18751
rect 543547 18687 543599 18693
rect 543555 18683 543591 18687
rect 543639 18667 543675 47920
rect 544808 47872 544844 59243
rect 543723 47836 544844 47872
rect 543631 18661 543683 18667
rect 543631 18603 543683 18609
rect 543639 18599 543675 18603
rect 543723 18583 543759 47836
rect 544892 47788 544928 59327
rect 561020 59271 561048 60454
rect 561260 60140 561288 60146
rect 561250 60134 561302 60140
rect 561502 60089 561538 60495
rect 561574 60187 561610 60540
rect 561646 60374 561682 60541
rect 561646 60346 561848 60374
rect 561250 60076 561302 60082
rect 561140 59852 561168 59856
rect 561128 59846 561180 59852
rect 561128 59788 561180 59794
rect 561140 59372 561168 59788
rect 561260 59442 561288 60076
rect 561700 59780 561728 59784
rect 561690 59774 561742 59780
rect 561690 59716 561742 59722
rect 561260 59414 561488 59442
rect 561140 59344 561368 59372
rect 561020 59243 561248 59271
rect 543807 47752 544928 47788
rect 543715 18577 543767 18583
rect 543715 18519 543767 18525
rect 543723 18515 543759 18519
rect 543807 18499 543843 47752
rect 555796 47465 556766 47742
rect 560962 47708 561014 47714
rect 560962 47650 561014 47656
rect 560722 47468 560774 47474
rect 560722 47410 560774 47416
rect 554946 46782 555918 47281
rect 546904 34216 547874 34482
rect 554946 34180 555916 34460
rect 558400 34014 559370 34549
rect 550056 33145 551028 33532
rect 554646 33409 555618 33968
rect 558128 28626 558136 28658
rect 559043 28626 559051 28658
rect 558128 27705 559051 28626
rect 546604 20228 547574 21098
rect 550056 20713 551026 21119
rect 546604 20108 546844 20228
rect 547192 20108 547574 20228
rect 554646 20214 555616 21084
rect 554646 20120 554920 20214
rect 554640 20108 554920 20120
rect 555294 20108 555616 20214
rect 558100 20099 559070 21082
rect 543799 18493 543851 18499
rect 543799 18435 543851 18441
rect 543807 18433 543843 18435
rect 560740 17838 560768 47410
rect 560844 47348 560896 47354
rect 560844 47290 560896 47296
rect 542752 17810 560768 17838
rect 542640 8538 542668 8556
rect 542622 8532 542674 8538
rect 542622 8474 542674 8480
rect 542528 8454 542556 8464
rect 542510 8448 542562 8454
rect 542510 8390 542562 8396
rect 542398 8364 542450 8370
rect 542398 8306 542450 8312
rect 542286 8280 542338 8288
rect 542286 8222 542338 8228
rect 542192 8202 542220 8204
rect 542174 8196 542226 8202
rect 542174 8138 542226 8144
rect 542080 8118 542108 8128
rect 542062 8112 542114 8118
rect 542062 8054 542114 8060
rect 541968 8034 541996 8042
rect 541950 8028 542002 8034
rect 541950 7970 542002 7976
rect 541856 7950 541884 7960
rect 541838 7944 541890 7950
rect 541838 7886 541890 7892
rect 541744 7866 541772 7868
rect 541726 7860 541778 7866
rect 541726 7802 541778 7808
rect 541632 7782 541660 7786
rect 541618 7776 541670 7782
rect 541618 7718 541670 7724
rect 541520 7698 541548 7712
rect 541510 7692 541562 7698
rect 541510 7634 541562 7640
rect 541408 7614 541436 7620
rect 541402 7608 541454 7614
rect 541402 7550 541454 7556
rect 541296 7530 541324 7538
rect 541290 7524 541342 7530
rect 541290 7466 541342 7472
rect 541184 7446 541212 7452
rect 541178 7440 541230 7446
rect 541178 7382 541230 7388
rect 541072 7362 541100 7366
rect 541066 7356 541118 7362
rect 541066 7298 541118 7304
rect 540960 7278 540988 7284
rect 540954 7272 541006 7278
rect 540954 7214 541006 7220
rect 540848 7194 540876 7198
rect 540840 7188 540892 7194
rect 540840 7130 540892 7136
rect 540736 7110 540764 7112
rect 540726 7104 540778 7110
rect 540726 7046 540778 7052
rect 540624 7026 540652 7034
rect 540612 7020 540664 7026
rect 540612 6962 540664 6968
rect 540512 6942 540540 6950
rect 540498 6936 540550 6942
rect 540498 6878 540550 6884
rect 540400 6858 540428 6862
rect 540384 6852 540436 6858
rect 540384 6794 540436 6800
rect 540400 0 540428 6794
rect 540512 0 540540 6878
rect 540624 0 540652 6962
rect 540736 0 540764 7046
rect 540848 0 540876 7130
rect 540960 0 540988 7214
rect 541072 0 541100 7298
rect 541184 0 541212 7382
rect 541296 0 541324 7466
rect 541408 0 541436 7550
rect 541520 0 541548 7634
rect 541632 0 541660 7718
rect 541744 0 541772 7802
rect 541856 0 541884 7886
rect 541968 0 541996 7970
rect 542080 0 542108 8054
rect 542192 0 542220 8138
rect 542304 0 542332 8222
rect 542416 0 542444 8306
rect 542528 0 542556 8390
rect 542640 0 542668 8474
rect 542752 0 542780 17810
rect 560860 17718 560888 47290
rect 542864 17690 560888 17718
rect 542864 0 542892 17690
rect 560980 17598 561008 47650
rect 561088 47594 561140 47600
rect 561088 47536 561140 47542
rect 542976 17570 561008 17598
rect 542976 0 543004 17570
rect 561100 17478 561128 47536
rect 543088 17450 561128 17478
rect 543088 0 543116 17450
rect 561220 17358 561248 59243
rect 543424 17330 561248 17358
rect 543200 14758 543228 14762
rect 543188 14752 543240 14758
rect 543188 14694 543240 14700
rect 543200 0 543228 14694
rect 543300 5337 543352 5343
rect 543300 5279 543352 5285
rect 543312 0 543340 5279
rect 543424 0 543452 17330
rect 561340 17238 561368 59344
rect 544208 17210 561368 17238
rect 543984 14838 544012 14840
rect 543972 14832 544024 14838
rect 543972 14774 544024 14780
rect 543536 0 543564 10578
rect 543648 0 543676 10657
rect 543760 0 543788 10727
rect 543872 0 543900 10792
rect 543984 0 544012 14774
rect 544084 5251 544136 5257
rect 544084 5193 544136 5199
rect 544096 0 544124 5193
rect 544208 0 544236 17210
rect 561460 17118 561488 59414
rect 561580 48114 561608 48120
rect 561570 48108 561622 48114
rect 561570 48050 561622 48056
rect 544880 17090 561488 17118
rect 544656 14928 544684 14932
rect 544644 14922 544696 14928
rect 544644 14864 544696 14870
rect 544320 0 544348 10876
rect 544432 0 544460 10939
rect 544544 0 544572 11018
rect 544656 0 544684 14864
rect 544756 5167 544808 5173
rect 544756 5109 544808 5115
rect 544768 0 544796 5109
rect 544880 0 544908 17090
rect 561580 16998 561608 48050
rect 545664 16970 561608 16998
rect 545440 15012 545468 15014
rect 545428 15006 545480 15012
rect 545428 14948 545480 14954
rect 544992 0 545020 11095
rect 545104 0 545132 11162
rect 545216 0 545244 11239
rect 545328 0 545356 11320
rect 545440 0 545468 14948
rect 545540 5084 545592 5090
rect 545540 5026 545592 5032
rect 545552 0 545580 5026
rect 545664 0 545692 16970
rect 561700 16878 561728 59716
rect 546112 16850 561728 16878
rect 545776 0 545804 11392
rect 545888 0 545916 11465
rect 546000 0 546028 11541
rect 546112 0 546140 16850
rect 561820 16758 561848 60346
rect 561940 60234 561968 60238
rect 562697 60236 562759 60665
rect 564261 60236 564300 60665
rect 561926 60228 561978 60234
rect 561926 60170 561978 60176
rect 546448 16730 561848 16758
rect 546224 0 546252 11611
rect 546336 0 546364 11673
rect 546448 0 546476 16730
rect 561940 16638 561968 60170
rect 562697 60167 564300 60236
rect 562420 60152 562448 60162
rect 562408 60146 562460 60152
rect 562408 60088 562460 60094
rect 562060 60068 562088 60074
rect 562048 60062 562100 60068
rect 562048 60004 562100 60010
rect 546896 16610 561968 16638
rect 546560 0 546588 11762
rect 546672 0 546700 11824
rect 546784 0 546812 11907
rect 546896 0 546924 16610
rect 562060 16518 562088 60004
rect 562180 59708 562208 59714
rect 562168 59702 562220 59708
rect 562168 59644 562220 59650
rect 547344 16490 562088 16518
rect 547008 0 547036 11977
rect 547120 0 547148 12054
rect 547232 0 547260 12121
rect 547344 0 547372 16490
rect 562180 16398 562208 59644
rect 562300 48034 562328 48038
rect 562288 48028 562340 48034
rect 562288 47970 562340 47976
rect 547680 16370 562208 16398
rect 547456 0 547484 12209
rect 547568 0 547596 12281
rect 547680 0 547708 16370
rect 562300 16278 562328 47970
rect 548128 16250 562328 16278
rect 547792 0 547820 12343
rect 547904 0 547932 12417
rect 548016 0 548044 12494
rect 548128 0 548156 16250
rect 562420 16158 562448 60088
rect 562660 59996 562688 60002
rect 562646 59990 562698 59996
rect 562646 59932 562698 59938
rect 562540 59636 562568 59640
rect 562528 59630 562580 59636
rect 562528 59572 562580 59578
rect 550256 16130 562448 16158
rect 550144 15176 550172 15180
rect 550132 15170 550184 15176
rect 550132 15112 550184 15118
rect 549808 15098 549836 15104
rect 549796 15092 549848 15098
rect 549796 15034 549848 15040
rect 548240 0 548268 12566
rect 548352 0 548380 12645
rect 548464 0 548492 12719
rect 548576 0 548604 12785
rect 548688 0 548716 12859
rect 548800 0 548828 12951
rect 548912 0 548940 13026
rect 549024 0 549052 13098
rect 549136 0 549164 13159
rect 549248 0 549276 13238
rect 549348 5001 549400 5007
rect 549348 4943 549400 4949
rect 549360 0 549388 4943
rect 549460 4917 549512 4923
rect 549460 4859 549512 4865
rect 549472 0 549500 4859
rect 549572 4834 549624 4840
rect 549572 4776 549624 4782
rect 549584 0 549612 4776
rect 549684 4749 549736 4755
rect 549684 4691 549736 4697
rect 549696 0 549724 4691
rect 549808 0 549836 15034
rect 549908 4666 549960 4672
rect 549908 4608 549960 4614
rect 549920 0 549948 4608
rect 550020 4580 550072 4586
rect 550020 4522 550072 4528
rect 550032 0 550060 4522
rect 550144 0 550172 15112
rect 550256 0 550284 16130
rect 562540 16038 562568 59572
rect 551264 16010 562568 16038
rect 551152 15428 551180 15432
rect 551140 15422 551192 15428
rect 551140 15364 551192 15370
rect 551040 15346 551068 15348
rect 551028 15340 551080 15346
rect 551028 15282 551080 15288
rect 550704 15260 550732 15264
rect 550692 15254 550744 15260
rect 550692 15196 550744 15202
rect 550368 0 550396 13332
rect 550480 0 550508 13332
rect 550592 0 550620 13424
rect 550704 0 550732 15196
rect 550804 4497 550856 4503
rect 550804 4439 550856 4445
rect 550816 0 550844 4439
rect 550916 4414 550968 4420
rect 550916 4356 550968 4362
rect 550928 0 550956 4356
rect 551040 0 551068 15282
rect 551152 0 551180 15364
rect 551264 0 551292 16010
rect 552608 15918 552636 15958
rect 562660 15918 562688 59932
rect 564812 59924 564840 59932
rect 564801 59918 564854 59924
rect 564853 59866 564854 59918
rect 564801 59860 564854 59866
rect 562780 47954 562808 47962
rect 562770 47948 562822 47954
rect 562770 47890 562822 47896
rect 552608 15890 562688 15918
rect 552484 15592 552536 15598
rect 552484 15534 552536 15540
rect 552160 15510 552188 15522
rect 552148 15504 552200 15510
rect 552148 15446 552200 15452
rect 551376 0 551404 13510
rect 551488 0 551516 13510
rect 551600 0 551628 13654
rect 551700 4327 551752 4333
rect 551700 4269 551752 4275
rect 551712 0 551740 4269
rect 551812 4244 551864 4250
rect 551812 4186 551864 4192
rect 551824 0 551852 4186
rect 551924 4160 551976 4166
rect 551924 4102 551976 4108
rect 551936 0 551964 4102
rect 552036 4076 552088 4082
rect 552036 4018 552088 4024
rect 552048 0 552076 4018
rect 552160 0 552188 15446
rect 552260 3993 552312 3999
rect 552260 3935 552312 3941
rect 552272 0 552300 3935
rect 552372 3908 552424 3914
rect 552372 3850 552424 3856
rect 552384 0 552412 3850
rect 552496 0 552524 15534
rect 552608 0 552636 15890
rect 553380 15842 553432 15848
rect 562780 15798 562808 47890
rect 562900 47874 562928 47882
rect 562886 47868 562938 47874
rect 562886 47810 562938 47816
rect 553380 15784 553432 15790
rect 553268 15756 553320 15762
rect 553268 15698 553320 15704
rect 552932 15674 552984 15680
rect 552932 15616 552984 15622
rect 552720 0 552748 13750
rect 552832 0 552860 13750
rect 552944 0 552972 15616
rect 553044 3824 553096 3830
rect 553044 3766 553096 3772
rect 553056 0 553084 3766
rect 553156 3742 553208 3748
rect 553156 3684 553208 3690
rect 553168 0 553196 3684
rect 553280 0 553308 15698
rect 553392 0 553420 15784
rect 553504 15770 562808 15798
rect 553504 0 553532 15770
rect 562900 15678 562928 47810
rect 554624 15650 562928 15678
rect 553616 0 553644 13942
rect 553728 0 553756 14010
rect 553840 0 553868 14080
rect 553940 3656 553992 3662
rect 553940 3598 553992 3604
rect 553952 0 553980 3598
rect 554052 3572 554104 3578
rect 554052 3514 554104 3520
rect 554064 0 554092 3514
rect 554164 3488 554216 3494
rect 554164 3430 554216 3436
rect 554176 0 554204 3430
rect 554276 3404 554328 3410
rect 554276 3346 554328 3352
rect 554288 0 554316 3346
rect 554388 3321 554440 3327
rect 554388 3263 554440 3269
rect 554400 0 554428 3263
rect 554500 3237 554552 3243
rect 554500 3179 554552 3185
rect 554512 0 554540 3179
rect 554624 0 554652 15650
rect 563020 15558 563048 58264
rect 555520 15530 563048 15558
rect 554736 0 554764 14164
rect 554848 0 554876 14228
rect 554948 3154 555000 3160
rect 554948 3096 555000 3102
rect 554960 0 554988 3096
rect 555060 3068 555112 3074
rect 555060 3010 555112 3016
rect 555072 0 555100 3010
rect 555184 0 555212 14296
rect 555296 0 555324 14362
rect 555408 0 555436 14448
rect 555520 0 555548 15530
rect 563132 15446 563160 58146
rect 555632 15418 563160 15446
rect 555632 0 555660 15418
rect 563244 15334 563272 58014
rect 555744 15306 563272 15334
rect 555744 0 555772 15306
rect 563356 15222 563384 57892
rect 555856 15194 563384 15222
rect 555856 0 555884 15194
rect 563468 15110 563496 57770
rect 555968 15082 563496 15110
rect 555968 0 555996 15082
rect 563580 14998 563608 57654
rect 556080 14970 563608 14998
rect 556080 0 556108 14970
rect 563692 14886 563720 57532
rect 556192 14858 563720 14886
rect 556192 0 556220 14858
rect 563804 14774 563832 57418
rect 556304 14746 563832 14774
rect 556304 0 556332 14746
rect 563916 14662 563944 57300
rect 556416 14634 563944 14662
rect 556416 0 556444 14634
rect 564028 14550 564056 57180
rect 556528 14522 564056 14550
rect 556528 0 556556 14522
rect 564140 14438 564168 57058
rect 556640 14410 564168 14438
rect 556640 0 556668 14410
rect 564252 14326 564280 56942
rect 556752 14298 564280 14326
rect 556752 0 556780 14298
rect 564364 14214 564392 56824
rect 556864 14186 564392 14214
rect 556864 0 556892 14186
rect 564476 14102 564504 56710
rect 556976 14074 564504 14102
rect 556976 0 557004 14074
rect 564588 13990 564616 56594
rect 557088 13962 564616 13990
rect 557088 0 557116 13962
rect 564700 13878 564728 56474
rect 557200 13850 564728 13878
rect 557200 0 557228 13850
rect 564812 13748 564840 59860
rect 565173 58968 566648 58997
rect 565173 58543 565210 58968
rect 566611 58543 566648 58968
rect 565173 58514 566648 58543
rect 566822 56241 566850 79865
rect 568948 79781 568976 88814
rect 569060 88758 569088 88768
rect 569048 88752 569100 88758
rect 569048 88694 569100 88700
rect 557312 13720 564840 13748
rect 565036 56213 566850 56241
rect 566934 79753 568976 79781
rect 557312 -20 557340 13720
rect 565036 13542 565064 56213
rect 566934 56129 566962 79753
rect 569060 79669 569088 88694
rect 569172 88624 569200 88630
rect 569160 88618 569212 88624
rect 569160 88560 569212 88566
rect 557536 13514 565064 13542
rect 565148 56101 566962 56129
rect 567046 79641 569088 79669
rect 557536 0 557564 13514
rect 565148 13430 565176 56101
rect 567046 56017 567074 79641
rect 569172 79557 569200 88560
rect 569284 83080 569312 83086
rect 569272 83074 569324 83080
rect 569272 83016 569324 83022
rect 557648 13402 565176 13430
rect 565260 55989 567074 56017
rect 567158 79529 569200 79557
rect 557648 0 557676 13402
rect 565260 13318 565288 55989
rect 567158 55905 567186 79529
rect 569284 79445 569312 83016
rect 569396 82962 569424 82968
rect 569384 82956 569436 82962
rect 569384 82898 569436 82904
rect 557760 13290 565288 13318
rect 565372 55877 567186 55905
rect 567270 79417 569312 79445
rect 557760 0 557788 13290
rect 565372 13206 565400 55877
rect 567270 55793 567298 79417
rect 569396 79333 569424 82898
rect 569508 82842 569536 82854
rect 569496 82836 569548 82842
rect 569496 82778 569548 82784
rect 557872 13178 565400 13206
rect 565484 55765 567298 55793
rect 567382 79305 569424 79333
rect 557872 0 557900 13178
rect 565484 13094 565512 55765
rect 567382 55681 567410 79305
rect 569508 79221 569536 82778
rect 569620 82728 569648 82734
rect 569608 82722 569660 82728
rect 569608 82664 569660 82670
rect 557984 13066 565512 13094
rect 565596 55653 567410 55681
rect 567494 79193 569536 79221
rect 557984 0 558012 13066
rect 565596 12982 565624 55653
rect 567494 55569 567522 79193
rect 569620 79109 569648 82664
rect 558096 12954 565624 12982
rect 565708 55541 567522 55569
rect 567606 79081 569648 79109
rect 558096 0 558124 12954
rect 565708 12870 565736 55541
rect 567606 55457 567634 79081
rect 569728 78962 569768 110382
rect 567728 78922 569768 78962
rect 567728 58192 567768 78922
rect 569848 78842 569888 110508
rect 567848 78802 569888 78842
rect 567848 58080 567888 78802
rect 569968 78722 570008 110612
rect 567968 78682 570008 78722
rect 567968 57964 568008 78682
rect 570088 78602 570128 110732
rect 568088 78562 570128 78602
rect 568088 57840 568128 78562
rect 570208 78482 570248 110852
rect 568208 78442 570248 78482
rect 568208 57722 568248 78442
rect 570328 78362 570368 110972
rect 568328 78322 570368 78362
rect 568328 57608 568368 78322
rect 570448 78242 570488 111092
rect 568448 78202 570488 78242
rect 568448 57488 568488 78202
rect 570568 78122 570608 111212
rect 568568 78082 570608 78122
rect 568568 57366 568608 78082
rect 570688 78002 570728 111332
rect 568688 77962 570728 78002
rect 568688 57254 568728 77962
rect 570808 77882 570848 111452
rect 568808 77842 570848 77882
rect 568808 57122 568848 77842
rect 570928 77762 570968 111572
rect 568928 77722 570968 77762
rect 568928 57004 568968 77722
rect 571048 77642 571088 111692
rect 569048 77602 571088 77642
rect 569048 56880 569088 77602
rect 571168 77522 571208 111812
rect 569168 77482 571208 77522
rect 569168 56770 569208 77482
rect 571288 77402 571328 111932
rect 569288 77362 571328 77402
rect 569288 56650 569328 77362
rect 571408 77282 571448 112052
rect 569408 77242 571448 77282
rect 569408 56528 569448 77242
rect 571528 77162 571568 112172
rect 569528 77122 571568 77162
rect 569528 56410 569568 77122
rect 558208 12842 565736 12870
rect 565820 55429 567634 55457
rect 558208 0 558236 12842
rect 565820 12758 565848 55429
rect 568620 54676 568648 54694
rect 568608 54670 568660 54676
rect 568608 54612 568660 54618
rect 567724 54426 567752 54432
rect 567712 54420 567764 54426
rect 567712 54362 567764 54368
rect 567500 48768 567528 48778
rect 567488 48762 567540 48768
rect 567488 48704 567540 48710
rect 567276 48528 567304 48534
rect 567264 48522 567316 48528
rect 567264 48464 567316 48470
rect 567052 41442 567080 41450
rect 567040 41436 567092 41442
rect 567040 41378 567092 41384
rect 566828 41188 566856 41194
rect 566816 41182 566868 41188
rect 566816 41124 566868 41130
rect 566604 35536 566632 35544
rect 566592 35530 566644 35536
rect 566592 35472 566644 35478
rect 566380 35302 566408 35308
rect 566368 35296 566420 35302
rect 566368 35238 566420 35244
rect 566156 28044 566184 28052
rect 566144 28038 566196 28044
rect 566144 27980 566196 27986
rect 565932 27822 565960 27828
rect 565920 27816 565972 27822
rect 565920 27758 565972 27764
rect 558320 12730 565848 12758
rect 558320 0 558348 12730
rect 565932 12646 565960 27758
rect 566044 27692 566072 27700
rect 566032 27686 566084 27692
rect 566032 27628 566084 27634
rect 558432 12618 565960 12646
rect 558432 0 558460 12618
rect 566044 12534 566072 27628
rect 558544 12506 566072 12534
rect 558544 0 558572 12506
rect 566156 12422 566184 27980
rect 566268 27936 566296 27944
rect 566256 27930 566308 27936
rect 566256 27872 566308 27878
rect 558656 12394 566184 12422
rect 558656 0 558684 12394
rect 566268 12310 566296 27872
rect 558768 12282 566296 12310
rect 558768 0 558796 12282
rect 566380 12198 566408 35238
rect 566492 35162 566520 35172
rect 566480 35156 566532 35162
rect 566480 35098 566532 35104
rect 558880 12170 566408 12198
rect 558880 0 558908 12170
rect 566492 12086 566520 35098
rect 558992 12058 566520 12086
rect 558992 0 559020 12058
rect 566604 11974 566632 35472
rect 566716 35408 566744 35424
rect 566704 35402 566756 35408
rect 566704 35344 566756 35350
rect 559104 11946 566632 11974
rect 559104 0 559132 11946
rect 566716 11862 566744 35344
rect 559216 11834 566744 11862
rect 559216 0 559244 11834
rect 566828 11750 566856 41124
rect 566940 41084 566968 41092
rect 566928 41078 566980 41084
rect 566928 41020 566980 41026
rect 559328 11722 566856 11750
rect 559328 0 559356 11722
rect 566940 11638 566968 41020
rect 559440 11610 566968 11638
rect 559440 0 559468 11610
rect 567052 11526 567080 41378
rect 567164 41320 567192 41330
rect 567152 41314 567204 41320
rect 567152 41256 567204 41262
rect 559552 11498 567080 11526
rect 559552 0 559580 11498
rect 567164 11414 567192 41256
rect 559664 11386 567192 11414
rect 559664 0 559692 11386
rect 567276 11302 567304 48464
rect 567388 48404 567416 48410
rect 567376 48398 567428 48404
rect 567376 48340 567428 48346
rect 559776 11274 567304 11302
rect 559776 0 559804 11274
rect 567388 11190 567416 48340
rect 559888 11162 567416 11190
rect 559888 0 559916 11162
rect 567500 11078 567528 48704
rect 567612 48654 567640 48660
rect 567600 48648 567652 48654
rect 567600 48590 567652 48596
rect 560000 11050 567528 11078
rect 560000 0 560028 11050
rect 567612 10966 567640 48590
rect 560112 10938 567640 10966
rect 560112 0 560140 10938
rect 567724 10854 567752 54362
rect 567836 54318 567864 54328
rect 567824 54312 567876 54318
rect 567824 54254 567876 54260
rect 560224 10826 567752 10854
rect 560224 0 560252 10826
rect 567836 10742 567864 54254
rect 567948 47182 567976 47196
rect 567936 47176 567988 47182
rect 567936 47118 567988 47124
rect 560336 10714 567864 10742
rect 560336 0 560364 10714
rect 567948 10630 567976 47118
rect 568060 47058 568088 47074
rect 568048 47052 568100 47058
rect 568048 46994 568100 47000
rect 560448 10602 567976 10630
rect 560448 0 560476 10602
rect 568060 10518 568088 46994
rect 568396 34762 568424 34772
rect 568384 34756 568436 34762
rect 568384 34698 568436 34704
rect 568172 33526 568200 33534
rect 568160 33520 568212 33526
rect 568160 33462 568212 33468
rect 560560 10490 568088 10518
rect 560560 0 560588 10490
rect 568172 10406 568200 33462
rect 568284 33432 568312 33442
rect 568272 33426 568324 33432
rect 568272 33368 568324 33374
rect 560672 10378 568200 10406
rect 560672 0 560700 10378
rect 568284 10294 568312 33368
rect 560784 10266 568312 10294
rect 560784 0 560812 10266
rect 568396 10182 568424 34698
rect 568508 34618 568536 34630
rect 568496 34612 568548 34618
rect 568496 34554 568548 34560
rect 560896 10154 568424 10182
rect 560896 0 560924 10154
rect 568508 10070 568536 34554
rect 561008 10042 568536 10070
rect 561008 0 561036 10042
rect 568620 9958 568648 54612
rect 568732 54556 568760 54574
rect 568724 54550 568776 54556
rect 568724 54492 568776 54498
rect 561120 9930 568648 9958
rect 561120 0 561148 9930
rect 568732 9846 568760 54492
rect 569280 22144 569332 22150
rect 569280 22086 569332 22092
rect 568832 21890 568884 21896
rect 568832 21832 568884 21838
rect 561232 9818 568760 9846
rect 561232 0 561260 9818
rect 568844 9734 568872 21832
rect 568944 21788 568996 21794
rect 568944 21730 568996 21736
rect 561344 9706 568872 9734
rect 561344 0 561372 9706
rect 568956 9622 568984 21730
rect 569056 21670 569108 21676
rect 569056 21612 569108 21618
rect 561456 9594 568984 9622
rect 561456 0 561484 9594
rect 569068 9510 569096 21612
rect 569168 21562 569220 21568
rect 569168 21504 569220 21510
rect 561568 9482 569096 9510
rect 561568 0 561596 9482
rect 569180 9398 569208 21504
rect 561680 9370 569208 9398
rect 561680 0 561708 9370
rect 569292 9286 569320 22086
rect 569392 22022 569444 22028
rect 569392 21964 569444 21970
rect 561792 9258 569320 9286
rect 561792 0 561820 9258
rect 569404 9174 569432 21964
rect 569930 18824 570058 66978
rect 570246 9500 570374 64318
rect 570562 18824 570690 66978
rect 571194 18824 571322 66978
rect 561904 9146 569432 9174
rect 561904 0 561932 9146
rect 571510 8406 571638 63273
rect 571826 18824 571954 66978
rect 572142 8016 572270 62795
rect 572458 18824 572586 66978
<< via2 >>
rect 2511 64731 5983 65223
rect 154585 90232 156040 90355
rect 154673 88696 156003 88824
rect 47304 80913 47726 81226
rect 47304 79683 47726 79996
rect 81705 49721 81761 49777
rect 81620 49041 81676 49097
rect 81540 47681 81596 47737
rect 81451 47001 81507 47057
rect 81368 45641 81424 45697
rect 81285 41854 81341 41910
rect 81200 41504 81256 41560
rect 81116 41196 81172 41252
rect 81032 39115 81088 39171
rect 80946 38520 81002 38576
rect 160460 80742 160761 82089
rect 160996 80732 161307 81841
rect 193329 81115 193632 81893
rect 193852 81115 194157 82259
rect 198858 90469 200372 90609
rect 198845 88930 200359 89070
rect 84783 58525 84916 59287
rect 84782 50906 84925 51474
rect 84838 47335 84898 47395
rect 84836 47098 84896 47158
rect 84836 46587 84896 46647
rect 84806 39518 84866 39578
rect 84810 39178 84870 39238
rect 84806 38966 84866 39026
rect 183998 59273 185192 59797
rect 189798 58319 190768 58513
rect 182438 52513 183994 52696
rect 191120 54832 192099 55017
rect 186566 52384 187774 52604
rect 134394 47905 134530 48217
rect 186599 34181 188523 34827
rect 175103 31064 176317 31631
rect 90573 10985 90888 12520
rect 91116 10993 91423 11779
rect 123624 10977 123927 11829
rect 124147 10975 124449 12624
rect 175090 29146 176304 29713
rect 186663 28312 188472 28962
rect 244169 34357 246537 34975
rect 232705 31208 234494 31763
rect 232969 29312 234511 29867
rect 244399 28490 247152 29128
rect 257258 24982 257372 26004
rect 388908 90725 390258 90856
rect 388995 89177 390345 89308
rect 394851 80687 395147 82606
rect 395370 80671 395671 81462
rect 434187 90780 435612 90895
rect 434639 89231 435961 89367
rect 427385 80611 427699 81409
rect 427915 80638 428234 82532
rect 509759 83681 510920 83844
rect 509771 82541 510932 82704
rect 550814 82332 551597 82652
rect 294545 16433 295010 19081
rect 352180 58638 353960 59225
rect 341063 17816 341153 17906
rect 385274 43242 386087 43716
rect 384078 41169 385891 41614
rect 367625 40205 367732 40312
rect 543189 79844 544669 80189
rect 406725 59616 407761 59916
rect 403905 46006 404057 46464
rect 404206 46000 404358 46458
rect 421070 51773 421767 51919
rect 421046 48341 421743 48487
rect 420803 47023 421743 47148
rect 420789 46034 421670 46173
rect 384400 39126 385734 39680
rect 393779 32474 394848 32731
rect 430108 31573 430715 31890
rect 446720 44838 446789 45172
rect 446880 44838 446949 45172
rect 447040 44838 447109 45172
rect 447200 44838 447269 45172
rect 447360 44838 447429 45172
rect 447520 44838 447589 45172
rect 447680 44838 447749 45172
rect 447840 44838 447909 45172
rect 451596 44841 451665 45175
rect 451756 44841 451825 45175
rect 451916 44841 451985 45175
rect 452076 44841 452145 45175
rect 452236 44841 452305 45175
rect 452396 44841 452465 45175
rect 452556 44841 452625 45175
rect 452716 44841 452785 45175
rect 452125 41808 459416 42875
rect 473111 41785 480402 42852
rect 482109 44289 482416 44396
rect 392065 28615 392969 29084
rect 431923 21785 438850 22602
rect 464430 21538 464574 21999
rect 464722 21537 464866 21998
rect 465027 21536 465171 21997
rect 465360 21540 465504 22001
rect 467428 21539 467613 22000
rect 473177 21637 478353 22662
rect 367625 19589 367732 19696
rect 562759 60236 564261 60665
rect 565210 58543 566611 58968
<< metal3 >>
rect 80700 114450 103216 114650
rect 265777 114560 283501 114863
rect 283998 114549 289035 114862
rect 312386 114514 362012 114714
rect 504862 114556 528012 114756
rect 56808 114050 102344 114250
rect 222818 114192 280622 114392
rect 284814 114176 297212 114376
rect 491473 114284 503784 114518
rect 314180 114028 386012 114228
rect 32788 113650 91142 113850
rect 198756 113792 278940 113992
rect 504862 113956 505062 114556
rect 554128 114528 569900 114728
rect 551250 114198 552076 114258
rect 505803 113998 552076 114198
rect 551250 113958 552076 113998
rect 285636 113754 298012 113954
rect 327454 113646 410012 113846
rect 492728 113756 505062 113956
rect 554128 113730 554328 114528
rect 8826 113250 88968 113450
rect 174750 113392 265944 113592
rect 507025 113530 554328 113730
rect 329066 113210 434012 113410
rect 150802 112992 264646 113192
rect 508564 113116 570504 113244
rect 508564 112844 508692 113116
rect 8200 112716 508692 112844
rect 508910 112770 552022 112970
rect 508910 112570 509110 112770
rect 13588 112370 509110 112570
rect 509288 112494 552022 112622
rect 509288 112222 509416 112494
rect 13059 112094 509416 112222
rect 13125 111748 492606 111948
rect 13059 111472 492616 111600
rect 43901 111126 490988 111326
rect 12558 110850 490991 110978
rect 12558 110504 330924 110704
rect 12558 110228 506648 110356
rect 43433 109882 506648 110082
rect 508032 110004 511450 110014
rect 42797 109606 506648 109734
rect 508032 109535 508087 110004
rect 508795 109535 511450 110004
rect 508032 109514 511450 109535
rect 42812 109260 305222 109460
rect 42797 108984 305498 109112
rect 14317 107874 14847 108065
rect 14628 107865 14847 107874
rect 43403 107865 43815 108065
rect 90983 107522 91917 107808
rect 43619 107232 49336 107258
rect 43619 106779 43650 107232
rect 44525 106779 49336 107232
rect 43619 106758 49336 106779
rect 90983 105647 91269 107522
rect 283988 107382 288383 108358
rect 509033 108138 509653 108161
rect 509033 107636 509061 108138
rect 509627 108052 509653 108138
rect 509627 107782 511220 108052
rect 509627 107636 509653 107782
rect 509033 107611 509653 107636
rect 465217 106993 470598 107066
rect 233423 106448 239117 106546
rect 44897 105596 55023 105624
rect 44897 105047 44952 105596
rect 45825 105047 55023 105596
rect 44897 105026 55023 105047
rect 3326 102336 17708 102476
rect 13939 101999 14788 102199
rect 43387 101999 44419 102199
rect 4510 101726 22530 101866
rect 5686 101426 27360 101566
rect 2716 96480 32214 96620
rect 13433 96133 14788 96333
rect 43403 96133 44863 96333
rect 3892 95860 37066 96000
rect 5080 95560 41850 95700
rect 88338 92968 88688 93180
rect 174133 105837 176168 106058
rect 178513 105818 180543 106039
rect 233423 104915 234448 106448
rect 239019 104915 239117 106448
rect 233423 104817 239117 104915
rect 158151 96762 158956 96936
rect 195674 96747 196527 96921
rect 197181 95328 200098 95471
rect 154914 95068 157831 95211
rect 197787 94029 199634 94189
rect 155378 93769 157225 93929
rect 198391 92552 199997 92707
rect 155015 92292 156621 92447
rect 198816 90609 200405 90631
rect 198816 90469 198858 90609
rect 200372 90469 200405 90609
rect 198816 90451 200405 90469
rect 154532 90355 156082 90383
rect 5398 90038 28128 90252
rect 154532 90232 154585 90355
rect 156040 90232 156082 90355
rect 154532 90196 156082 90232
rect 5406 89464 20064 89678
rect 24668 89438 32833 89556
rect 16642 89042 32417 89168
rect 198814 89070 200403 89092
rect 198814 88930 198845 89070
rect 200359 88930 200403 89070
rect 198814 88912 200403 88930
rect 154634 88824 156048 88857
rect 154634 88696 154673 88824
rect 156003 88696 156048 88824
rect 154634 88671 156048 88696
rect 175449 88184 176238 88421
rect 178425 88164 179168 88401
rect 230261 85990 236699 86144
rect 230261 84812 230496 85990
rect 232362 84812 236699 85990
rect 230261 84632 236699 84812
rect 28033 84482 30615 84506
rect 28033 84214 28061 84482
rect 30580 84214 30615 84482
rect 28033 84191 30615 84214
rect 142669 82275 143743 82289
rect 142669 82140 142694 82275
rect 143519 82140 143743 82275
rect 142669 82110 143743 82140
rect 46156 81226 47751 81250
rect 46156 81190 47304 81226
rect 46156 80934 46174 81190
rect 46578 80934 47304 81190
rect 46156 80913 47304 80934
rect 47726 80913 47751 81226
rect 193813 82259 194192 82310
rect 160429 82089 160805 82143
rect 46156 80877 47751 80913
rect 44884 80778 49034 80796
rect 44884 80162 44940 80778
rect 45820 80162 49034 80778
rect 141492 80790 143708 80812
rect 141492 80655 141515 80790
rect 142340 80655 143708 80790
rect 160429 80742 160460 82089
rect 160761 80742 160805 82089
rect 193282 81893 193664 81934
rect 160429 80685 160805 80742
rect 160959 81841 161338 81881
rect 160959 80732 160996 81841
rect 161307 80732 161338 81841
rect 193282 81115 193329 81893
rect 193632 81115 193664 81893
rect 193282 81070 193664 81115
rect 193813 81115 193852 82259
rect 194157 81115 194192 82259
rect 211618 82253 215765 82425
rect 193813 81076 194192 81115
rect 211723 80936 215870 80949
rect 211723 80792 212513 80936
rect 213299 80792 215870 80936
rect 211723 80777 215870 80792
rect 211728 80769 213351 80777
rect 160959 80688 161338 80732
rect 141492 80633 143708 80655
rect 44884 80138 49034 80162
rect 198839 80135 199494 80147
rect 46826 79996 47751 80020
rect 46826 79960 47304 79996
rect 46826 79704 46844 79960
rect 47248 79704 47304 79960
rect 46826 79683 47304 79704
rect 47726 79683 47751 79996
rect 140419 80003 144108 80011
rect 140419 79863 140440 80003
rect 141141 79863 144108 80003
rect 140419 79847 144108 79863
rect 156806 79788 176224 80118
rect 178410 79788 198555 80118
rect 198839 79994 198863 80135
rect 199411 79994 199494 80135
rect 198839 79983 199494 79994
rect 211784 79975 215875 80146
rect 46826 79647 47751 79683
rect 139542 79442 144053 79454
rect 139542 79294 139559 79442
rect 140240 79294 144053 79442
rect 211784 79428 215875 79599
rect 139542 79280 144053 79294
rect 43572 79042 48844 79064
rect 43572 78584 43650 79042
rect 44534 78584 48844 79042
rect 43572 78564 48844 78584
rect 88973 78384 139937 78510
rect 16638 77958 32059 78092
rect 88973 77803 89099 78384
rect 139811 78110 139937 78384
rect 139811 77984 228260 78110
rect 263960 78038 264120 98936
rect 265622 78438 265782 106756
rect 278694 78838 278854 106682
rect 283996 103926 288695 104902
rect 280308 79238 280468 98766
rect 285610 95906 294806 96870
rect 283171 91266 288384 92244
rect 283170 87822 288727 88800
rect 284804 79816 294723 80802
rect 312420 79638 312580 98656
rect 314226 80038 314386 106676
rect 314930 90760 315326 91866
rect 315958 91574 316354 91876
rect 315958 91499 320210 91574
rect 315958 91178 319886 91499
rect 314930 90714 319366 90760
rect 314930 90364 319004 90714
rect 318970 88765 319004 90364
rect 319323 88765 319366 90714
rect 318970 88686 319366 88765
rect 319814 88736 319886 91178
rect 320160 88736 320210 91499
rect 319814 88671 320210 88736
rect 327366 80438 327526 106924
rect 409871 105385 410368 105606
rect 412713 105325 413210 105546
rect 465217 105291 465393 106993
rect 467127 105291 470598 106993
rect 465217 105107 470598 105291
rect 329092 80838 329252 98766
rect 392633 96312 393330 96486
rect 429748 96252 430727 96426
rect 389284 95558 392201 95701
rect 432351 95588 435268 95731
rect 550760 95724 551233 95936
rect 559056 95095 573719 95102
rect 559056 94802 573665 95095
rect 389748 94259 391595 94419
rect 432957 94289 434804 94449
rect 567097 94280 573056 94580
rect 389385 92782 390991 92937
rect 433561 92812 435167 92967
rect 434140 90895 435650 90933
rect 388877 90856 390307 90889
rect 388877 90725 388908 90856
rect 390258 90725 390307 90856
rect 434140 90780 434187 90895
rect 435612 90780 435650 90895
rect 434140 90741 435650 90780
rect 388877 90694 390307 90725
rect 434605 89395 435575 89397
rect 434605 89367 436007 89395
rect 388959 89308 390389 89349
rect 388959 89177 388995 89308
rect 390345 89177 390389 89308
rect 434605 89231 434639 89367
rect 435961 89231 436007 89367
rect 434605 89197 436007 89231
rect 388959 89154 390389 89177
rect 409857 87734 410438 87971
rect 412625 87674 413206 87911
rect 469860 86252 475470 86361
rect 469860 84830 473636 86252
rect 475432 84830 475470 86252
rect 489058 85106 508003 85271
rect 469860 84752 475470 84830
rect 499925 84146 500259 84185
rect 329092 80698 360690 80838
rect 394813 82606 395187 82661
rect 394813 80687 394851 82606
rect 395147 80687 395187 82606
rect 427887 82532 428279 82593
rect 394813 80638 395187 80687
rect 395338 81462 395710 81521
rect 395338 80671 395370 81462
rect 395671 80671 395710 81462
rect 395338 80627 395710 80671
rect 427342 81409 427744 81455
rect 427342 80611 427385 81409
rect 427699 80611 427744 81409
rect 427342 80571 427744 80611
rect 427887 80638 427915 82532
rect 428234 80638 428279 82532
rect 499925 82893 499949 84146
rect 500235 83864 500259 84146
rect 500235 83844 510951 83864
rect 500235 83681 509759 83844
rect 510920 83681 510951 83844
rect 500235 83662 510951 83681
rect 500235 82893 500259 83662
rect 509039 83514 511612 83552
rect 499925 82858 500259 82893
rect 501123 83150 501449 83194
rect 501123 82721 501152 83150
rect 501121 82519 501152 82721
rect 448369 82306 454714 82485
rect 501123 81984 501152 82519
rect 501407 82721 501449 83150
rect 509039 82928 509068 83514
rect 509620 82928 511612 83514
rect 509039 82894 511612 82928
rect 545932 83115 546947 83136
rect 501407 82704 510960 82721
rect 501407 82541 509771 82704
rect 510932 82541 510960 82704
rect 501407 82519 510960 82541
rect 501407 81984 501449 82519
rect 545932 82338 545974 83115
rect 546865 82688 546947 83115
rect 550773 82688 551644 82693
rect 546865 82652 551644 82688
rect 546865 82338 550814 82652
rect 545932 82332 550814 82338
rect 551597 82332 551644 82652
rect 545932 82283 551644 82332
rect 550773 82281 551644 82283
rect 501123 81945 501449 81984
rect 508082 82112 517176 82133
rect 508082 81348 508114 82112
rect 508775 81348 517176 82112
rect 508082 81320 517176 81348
rect 551786 81172 551980 84464
rect 448330 80829 454708 81008
rect 546076 80978 551980 81172
rect 427887 80581 428279 80638
rect 327366 80298 360248 80438
rect 448349 80303 454713 80320
rect 448349 80161 450757 80303
rect 451373 80161 454713 80303
rect 448349 80144 454713 80161
rect 375477 80126 376522 80141
rect 314226 79898 359700 80038
rect 375477 79999 375497 80126
rect 376097 79999 376522 80126
rect 375477 79977 376522 79999
rect 312420 79500 359170 79638
rect 312632 79498 359170 79500
rect 374676 79563 376768 79584
rect 374676 79434 374700 79563
rect 375223 79434 376768 79563
rect 374676 79410 376768 79434
rect 389419 79388 410424 79718
rect 412610 79388 435608 79718
rect 448424 79631 454728 79650
rect 448424 79499 451681 79631
rect 452277 79499 454728 79631
rect 448424 79476 454728 79499
rect 280306 79098 358692 79238
rect 526669 78943 527019 80830
rect 543134 80189 544731 80250
rect 543134 79844 543189 80189
rect 544669 79844 544731 80189
rect 543134 79804 544731 79844
rect 278694 78698 358130 78838
rect 546076 78734 546270 80978
rect 552233 80873 552427 84405
rect 567525 83208 567556 83547
rect 557534 81670 564611 81864
rect 546564 80679 552427 80873
rect 265622 78298 357606 78438
rect 546564 78386 546758 80679
rect 556012 80575 556206 81660
rect 546983 80381 556206 80575
rect 370496 78188 370832 78193
rect 379948 78188 380284 78193
rect 384374 78188 384710 78193
rect 389000 78188 389336 78193
rect 398252 78188 398588 78193
rect 402878 78188 403214 78193
rect 407504 78188 407840 78193
rect 412130 78188 412466 78193
rect 416756 78188 417092 78193
rect 421382 78188 421718 78193
rect 426008 78188 426344 78193
rect 430934 78188 431270 78193
rect 435260 78188 435596 78193
rect 440056 78188 440392 78193
rect 444682 78188 445018 78193
rect 449138 78188 449474 78193
rect 453934 78188 454270 78193
rect 458590 78188 458926 78193
rect 463116 78188 463452 78193
rect 467842 78188 468178 78193
rect 472468 78188 472804 78193
rect 477094 78188 477430 78193
rect 481720 78188 482056 78193
rect 486346 78188 486682 78193
rect 490972 78188 491308 78193
rect 495598 78188 495934 78193
rect 499924 78188 500260 78193
rect 546983 78058 547177 80381
rect 557534 80237 557728 81670
rect 559056 81404 562360 81494
rect 559056 81194 572750 81404
rect 562060 81104 572750 81194
rect 567099 80440 572160 80740
rect 547553 80043 557728 80237
rect 263960 77900 357090 78038
rect 264180 77898 357090 77900
rect 54040 77633 89100 77803
rect 547553 77722 547747 80043
rect 103654 77498 356600 77638
rect 361084 77498 499162 77638
rect 102853 77098 356078 77238
rect 361582 77098 500562 77238
rect 6020 76724 20076 76938
rect 24642 76802 31672 76928
rect 6564 76286 28146 76500
rect 64591 74483 64824 76897
rect 89882 76698 355574 76838
rect 362098 76698 506390 76838
rect 74322 74786 74541 76492
rect 85120 74833 85339 76539
rect 89520 76298 355050 76438
rect 362584 76298 506810 76438
rect 151638 75918 554411 76046
rect 151638 75662 554406 75790
rect 147656 75406 560614 75534
rect 147656 75150 548174 75278
rect 147656 74894 558956 75022
rect 272850 74638 558956 74766
rect 439540 74635 440071 74638
rect 268608 74382 558956 74510
rect 268608 74126 549641 74254
rect 32714 73870 554542 73998
rect 384629 73742 385160 73743
rect 32714 73614 554470 73742
rect 32314 73358 554470 73486
rect 379475 73230 380006 73233
rect 32314 73102 548140 73230
rect 31908 72846 559235 72974
rect 31920 72590 559235 72718
rect 31450 72334 559235 72462
rect 207433 72206 207964 72208
rect 31522 72078 549967 72206
rect 35012 71822 556247 71950
rect 151820 71694 152351 71701
rect 35056 71566 556247 71694
rect 33934 71310 556247 71438
rect 147303 71182 147834 71192
rect 33930 71054 548174 71182
rect 33512 70798 560925 70926
rect 34183 70542 560925 70670
rect 32994 70286 560925 70414
rect 33719 70030 549960 70158
rect 33010 69774 549960 69902
rect 134791 69519 290687 69647
rect 346356 69518 506614 69646
rect 134505 69390 346544 69391
rect 134505 69263 504468 69390
rect 346356 69262 504468 69263
rect 193175 69007 290384 69135
rect 346847 69006 506622 69134
rect 3051 68750 556542 68878
rect 2722 68494 556542 68622
rect 3665 68238 556542 68366
rect 3316 67982 548162 68110
rect 4264 67726 560957 67854
rect 3912 67470 560957 67598
rect 4835 67214 551617 67342
rect 4486 66958 551608 67086
rect 5406 66702 544479 66830
rect 5090 66446 544479 66574
rect 6013 66190 544877 66318
rect 569876 66262 572606 66970
rect 5684 65934 544781 66062
rect 5993 65678 544781 65806
rect 130843 65422 476970 65550
rect 2423 65286 5727 65287
rect 10917 65286 14755 65344
rect 2423 65236 14755 65286
rect 2423 65223 7360 65236
rect 2423 64731 2511 65223
rect 5983 64731 7360 65223
rect 2423 64720 7360 64731
rect 8556 65195 14755 65236
rect 8556 64720 11043 65195
rect 2423 64662 11043 64720
rect 10917 64365 11043 64662
rect 14614 64365 14755 65195
rect 83261 65166 453924 65294
rect 83261 64910 453924 65038
rect 83261 64654 506398 64782
rect 191048 64398 506398 64526
rect 10917 64208 14755 64365
rect 191048 64142 570485 64270
rect 228994 63886 570436 64014
rect 4411 63630 571132 63758
rect 4537 63374 506364 63502
rect 4878 63118 571797 63246
rect 199473 62762 285736 62914
rect 290486 62862 571797 62990
rect 155749 62411 285226 62583
rect 52573 62033 284843 62179
rect 7666 61700 28318 61850
rect 48553 61749 155285 61802
rect 48553 61639 284444 61749
rect 155122 61586 284444 61639
rect 8092 61310 20270 61474
rect 23926 61182 35334 61304
rect 85322 61258 133776 61284
rect 15888 60720 34944 60854
rect 85322 60752 132948 61258
rect 133712 60752 133776 61258
rect 85322 60716 133776 60752
rect 284281 60759 284444 61586
rect 284697 61168 284843 62033
rect 285054 61583 285226 62411
rect 285584 61914 285736 62762
rect 289885 62606 572363 62734
rect 289885 62350 572363 62478
rect 289885 62094 572363 62222
rect 285584 61762 388552 61914
rect 405373 61829 422326 61941
rect 405373 61788 414932 61829
rect 285054 61411 387938 61583
rect 284697 61022 386403 61168
rect 85322 60442 85890 60716
rect 283176 60589 283522 60598
rect 284281 60596 392821 60759
rect 414838 60678 414932 61788
rect 415612 61788 422326 61829
rect 415612 60678 415704 61788
rect 484465 61752 526678 61892
rect 540363 61699 565771 62002
rect 540363 61368 540666 61699
rect 530062 61065 540666 61368
rect 541626 61245 556496 61548
rect 84763 59287 84944 59315
rect 85322 59301 86040 60442
rect 282170 60157 283556 60589
rect 414838 60575 415704 60678
rect 520440 60641 527376 61001
rect 319470 60232 319670 60265
rect 320310 60259 320510 60265
rect 283176 60150 283522 60157
rect 183932 59797 185250 59846
rect 84763 58525 84783 59287
rect 84916 58525 84944 59287
rect 28867 56270 30627 56309
rect 28867 56030 29923 56270
rect 30568 56030 30627 56270
rect 28867 55989 30627 56030
rect 84763 51474 84944 58525
rect 125998 59100 130836 59141
rect 125998 58260 130264 59100
rect 130786 58260 130836 59100
rect 183932 59273 183998 59797
rect 185192 59273 185250 59797
rect 320310 59977 320333 60259
rect 328850 60191 387150 60355
rect 183932 59224 185250 59273
rect 282266 58535 286272 59597
rect 319470 59512 319670 59950
rect 320310 59512 320510 59977
rect 328850 59508 328990 60191
rect 520440 60161 527926 60521
rect 405417 59916 406546 59943
rect 406677 59916 407807 59944
rect 405417 59616 405465 59916
rect 406501 59616 406725 59916
rect 407761 59616 407807 59916
rect 405417 59583 406546 59616
rect 406677 59583 407807 59616
rect 372242 59420 373515 59489
rect 352133 59225 363109 59265
rect 189741 58513 190803 58535
rect 189741 58319 189798 58513
rect 190768 58319 190803 58513
rect 189741 58275 190803 58319
rect 125998 58223 130836 58260
rect 125998 58028 129632 58063
rect 125998 57232 129052 58028
rect 129570 57232 129632 58028
rect 125998 57181 129632 57232
rect 125972 56982 130858 57021
rect 125972 56262 130252 56982
rect 130774 56262 130858 56982
rect 125972 56221 130858 56262
rect 125954 56024 132351 56061
rect 125954 55114 131492 56024
rect 132264 55114 132351 56024
rect 283982 55956 284338 55964
rect 282206 55524 284352 55956
rect 283982 55510 284338 55524
rect 343043 56049 343173 56392
rect 343555 56049 343685 56636
rect 344067 56049 344197 56950
rect 344579 56049 344709 57372
rect 345091 56049 345221 57661
rect 345603 56049 345733 58033
rect 346115 56049 346245 58224
rect 346627 56049 346757 58414
rect 347139 56049 347269 58819
rect 348675 56049 348805 57745
rect 349187 56049 349317 57968
rect 349699 56049 349829 58216
rect 350211 56049 350341 58464
rect 350723 56049 350853 58803
rect 351235 56049 351365 59183
rect 352133 58638 352180 59225
rect 353960 58638 363109 59225
rect 352133 58603 363109 58638
rect 372242 58463 372341 59420
rect 373424 58463 373515 59420
rect 372242 57783 373515 58463
rect 529537 58947 529936 59028
rect 529537 57678 529578 58947
rect 529863 57678 529936 58947
rect 529537 57604 529936 57678
rect 530062 55702 530362 61065
rect 535535 59924 535855 59965
rect 530546 58995 530945 59061
rect 530546 57726 530611 58995
rect 530896 57726 530945 58995
rect 535535 58682 535562 59924
rect 535808 58682 535855 59924
rect 535535 58641 535855 58682
rect 536449 59928 536769 59959
rect 536449 58686 536487 59928
rect 536733 58686 536769 59928
rect 536449 58635 536769 58686
rect 530546 57637 530945 57726
rect 476680 55177 484244 55277
rect 476771 55172 477576 55177
rect 125954 55061 132351 55114
rect 191072 55017 192134 55048
rect 125946 54865 133521 54901
rect 125946 54136 132702 54865
rect 133477 54136 133521 54865
rect 191072 54832 191120 55017
rect 192099 54832 192134 55017
rect 191072 54788 192134 54832
rect 125946 54101 133521 54136
rect 125966 53942 133548 53991
rect 125966 52870 132724 53942
rect 133492 52870 133548 53942
rect 125966 52816 133548 52870
rect 372625 52920 375352 52966
rect 182377 52696 184035 52741
rect 182377 52513 182438 52696
rect 183994 52513 184035 52696
rect 182377 52464 184035 52513
rect 186469 52604 187820 52655
rect 186469 52451 186566 52604
rect 186479 52384 186566 52451
rect 187774 52384 187820 52604
rect 372625 52579 374345 52920
rect 375302 52579 375352 52920
rect 372625 52543 375352 52579
rect 186479 52333 187820 52384
rect 421035 51919 421805 51943
rect 421035 51773 421070 51919
rect 421767 51773 421805 51919
rect 421035 51738 421805 51773
rect 84763 50906 84782 51474
rect 84925 50906 84944 51474
rect 284788 51323 285144 51334
rect 15870 49734 34484 49856
rect 81700 49779 81766 49782
rect 80861 49777 81766 49779
rect 80861 49721 81705 49777
rect 81761 49721 81766 49777
rect 80861 49719 81766 49721
rect 81700 49716 81766 49719
rect 84763 49685 84944 50906
rect 282344 50891 285200 51323
rect 284788 50880 285144 50891
rect 131454 50210 132317 50257
rect 131454 49685 131501 50210
rect 84763 49554 131501 49685
rect 132272 49554 132317 50210
rect 84763 49504 132317 49554
rect 364735 50211 364936 50237
rect 86014 49374 86645 49408
rect 81615 49099 81681 49102
rect 80833 49097 81696 49099
rect 80833 49041 81620 49097
rect 81676 49041 81696 49097
rect 80833 49039 81696 49041
rect 81615 49036 81681 49039
rect 8652 48600 20254 48726
rect 24842 48636 34107 48778
rect 86014 48708 86040 49374
rect 86615 48708 86645 49374
rect 364735 49357 364765 50211
rect 364915 49357 364936 50211
rect 364735 49322 364936 49357
rect 368252 49395 369247 49435
rect 368252 49227 368319 49395
rect 369200 49227 369247 49395
rect 368252 49193 369247 49227
rect 86014 48503 86645 48708
rect 421004 48487 421774 48515
rect 9204 48162 28318 48304
rect 134383 48217 134708 48292
rect 134383 47905 134394 48217
rect 134530 47905 134708 48217
rect 193308 48194 193530 48430
rect 421004 48341 421046 48487
rect 421743 48341 421774 48487
rect 421004 48310 421774 48341
rect 193308 48059 193540 48194
rect 193308 48004 193530 48059
rect 134383 47866 134708 47905
rect 9668 47700 28318 47850
rect 81535 47739 81601 47742
rect 80861 47737 81609 47739
rect 80861 47681 81540 47737
rect 81596 47681 81609 47737
rect 80861 47679 81609 47681
rect 81535 47676 81601 47679
rect 10187 47310 20270 47474
rect 84832 47395 84904 47426
rect 23976 47206 33657 47340
rect 84832 47335 84838 47395
rect 84898 47335 84904 47395
rect 84832 47163 84904 47335
rect 84831 47158 84904 47163
rect 84831 47098 84836 47158
rect 84896 47098 84904 47158
rect 84831 47093 84904 47098
rect 16832 46932 33350 47082
rect 81446 47059 81512 47062
rect 80847 47057 81521 47059
rect 80847 47001 81451 47057
rect 81507 47001 81521 47057
rect 80847 46999 81521 47001
rect 81446 46996 81512 46999
rect 84832 46652 84904 47093
rect 84831 46647 84904 46652
rect 84831 46587 84836 46647
rect 84896 46587 84904 46647
rect 84831 46582 84904 46587
rect 84832 46102 84904 46582
rect 125986 47192 130830 47223
rect 125986 46352 130254 47192
rect 130776 46352 130830 47192
rect 420754 47158 421778 47190
rect 420754 47148 421781 47158
rect 420754 47023 420803 47148
rect 421743 47023 421781 47148
rect 420754 46988 421781 47023
rect 285606 46690 285962 46702
rect 125986 46305 130830 46352
rect 282326 46258 285970 46690
rect 403880 46464 404079 46486
rect 285606 46248 285962 46258
rect 81359 46028 84904 46102
rect 125994 46104 129656 46145
rect 81363 45699 81429 45702
rect 80804 45697 81435 45699
rect 80804 45641 81368 45697
rect 81424 45641 81435 45697
rect 80804 45639 81435 45641
rect 81363 45636 81429 45639
rect 125994 45292 129052 46104
rect 129564 45292 129656 46104
rect 403880 46006 403905 46464
rect 404057 46006 404079 46464
rect 403880 45978 404079 46006
rect 404186 46458 404385 46486
rect 404186 46000 404206 46458
rect 404358 46000 404385 46458
rect 420747 46173 421736 46211
rect 420747 46034 420789 46173
rect 421670 46034 421736 46173
rect 420747 46003 421736 46034
rect 403756 45940 404086 45978
rect 125994 45263 129656 45292
rect 402878 45342 403415 45397
rect 125990 45079 130848 45103
rect 125990 44332 130246 45079
rect 130791 44332 130848 45079
rect 402878 44613 402922 45342
rect 403374 44767 403415 45342
rect 403756 44919 403806 45940
rect 404042 44919 404086 45940
rect 403756 44879 404086 44919
rect 403880 44875 404079 44879
rect 404186 44767 404385 46000
rect 446715 45172 446795 45218
rect 446715 44838 446720 45172
rect 446789 44838 446795 45172
rect 446715 44832 446795 44838
rect 446875 45172 446955 45218
rect 446875 44838 446880 45172
rect 446949 44838 446955 45172
rect 446875 44832 446955 44838
rect 447035 45172 447115 45218
rect 447035 44838 447040 45172
rect 447109 44838 447115 45172
rect 447035 44832 447115 44838
rect 447195 45172 447275 45218
rect 447195 44838 447200 45172
rect 447269 44838 447275 45172
rect 447195 44832 447275 44838
rect 447355 45172 447435 45218
rect 447355 44838 447360 45172
rect 447429 44838 447435 45172
rect 447355 44832 447435 44838
rect 447515 45172 447595 45218
rect 447515 44838 447520 45172
rect 447589 44838 447595 45172
rect 447515 44832 447595 44838
rect 447675 45172 447755 45218
rect 447675 44838 447680 45172
rect 447749 44838 447755 45172
rect 447675 44832 447755 44838
rect 447835 45172 447915 45218
rect 447835 44838 447840 45172
rect 447909 44838 447915 45172
rect 447835 44832 447915 44838
rect 451591 45175 451671 45192
rect 451591 44841 451596 45175
rect 451665 44841 451671 45175
rect 451591 44835 451671 44841
rect 451751 45175 451831 45192
rect 451751 44841 451756 45175
rect 451825 44841 451831 45175
rect 451751 44835 451831 44841
rect 451911 45175 451991 45192
rect 451911 44841 451916 45175
rect 451985 44841 451991 45175
rect 451911 44835 451991 44841
rect 452071 45175 452151 45192
rect 452071 44841 452076 45175
rect 452145 44841 452151 45175
rect 452071 44835 452151 44841
rect 452231 45175 452311 45192
rect 452231 44841 452236 45175
rect 452305 44841 452311 45175
rect 452231 44835 452311 44841
rect 452391 45175 452471 45192
rect 452391 44841 452396 45175
rect 452465 44841 452471 45175
rect 452391 44835 452471 44841
rect 452551 45175 452631 45192
rect 452551 44841 452556 45175
rect 452625 44841 452631 45175
rect 452551 44835 452631 44841
rect 452711 44841 452716 44966
rect 452785 44841 452791 44966
rect 452711 44835 452791 44841
rect 403374 44613 404385 44767
rect 421907 44652 436556 44757
rect 402878 44569 404385 44613
rect 402886 44568 404385 44569
rect 125990 44303 130848 44332
rect 367620 44430 390179 44547
rect 81338 44114 86044 44143
rect 81338 43170 81394 44114
rect 82156 43170 86044 44114
rect 81338 43143 86044 43170
rect 86014 42962 100674 42983
rect 28896 42289 30633 42313
rect 28896 42025 29917 42289
rect 30568 42025 30633 42289
rect 86014 42201 99918 42962
rect 100644 42201 100674 42962
rect 86014 42183 100674 42201
rect 28896 41993 30633 42025
rect 81280 41912 81346 41915
rect 80861 41910 81356 41912
rect 80861 41854 81285 41910
rect 81341 41854 81356 41910
rect 80861 41852 81356 41854
rect 81280 41849 81346 41852
rect 82769 41778 86024 41806
rect 81195 41562 81261 41565
rect 80835 41560 81270 41562
rect 80835 41504 81200 41560
rect 81256 41504 81270 41560
rect 80835 41502 81270 41504
rect 81195 41499 81261 41502
rect 81111 41254 81177 41257
rect 80849 41252 81181 41254
rect 80849 41196 81116 41252
rect 81172 41196 81181 41252
rect 80849 41194 81181 41196
rect 81111 41191 81177 41194
rect 82769 40922 82822 41778
rect 83516 40922 86024 41778
rect 82769 40888 86024 40922
rect 367620 40312 367737 44430
rect 390062 44401 390179 44430
rect 390062 44396 483829 44401
rect 390062 44289 482109 44396
rect 482416 44289 483829 44396
rect 390062 44284 483829 44289
rect 385241 43716 386119 43750
rect 484144 43739 484244 55177
rect 541626 54778 541929 61245
rect 550881 60812 565726 61112
rect 562697 60665 564307 60715
rect 544080 60176 556739 60304
rect 562697 60236 562759 60665
rect 564261 60236 564307 60665
rect 562697 60167 564307 60236
rect 544321 59827 548671 59955
rect 559248 59743 566350 60043
rect 565167 59030 567607 59053
rect 565167 58968 566623 59030
rect 565167 58543 565210 58968
rect 566611 58543 566623 58968
rect 565167 58523 566623 58543
rect 567534 58523 567607 59030
rect 565167 58502 567607 58523
rect 530096 49277 530406 52296
rect 541587 49280 541841 52255
rect 559248 51613 567490 51913
rect 530096 49023 540537 49277
rect 527662 47682 535758 47933
rect 530699 47402 539225 47409
rect 530696 47126 539225 47402
rect 540283 47090 540537 49023
rect 540862 49026 541841 49280
rect 540862 47090 541116 49026
rect 551206 48405 566922 48705
rect 543863 47551 548704 47679
rect 549336 47457 556775 47585
rect 549336 47390 549464 47457
rect 543593 47262 549464 47390
rect 549712 47124 555919 47252
rect 549712 47113 549840 47124
rect 543066 46985 549840 47113
rect 543317 46718 547871 46846
rect 550356 46579 568126 46879
rect 558397 44263 568752 44563
rect 385241 43242 385274 43716
rect 386087 43242 386119 43716
rect 482857 43639 484244 43739
rect 435475 43313 461616 43477
rect 385241 43211 386119 43242
rect 451969 42875 459639 43075
rect 451969 41808 452125 42875
rect 459416 41808 459639 42875
rect 461452 42849 461616 43313
rect 479068 43008 480580 43009
rect 472888 42852 480580 43008
rect 384012 41614 385956 41662
rect 384012 41169 384078 41614
rect 385891 41169 385956 41614
rect 451969 41608 459639 41808
rect 472888 41785 473111 42852
rect 480402 41785 480580 42852
rect 472888 41541 480580 41785
rect 384012 41112 385956 41169
rect 367620 40205 367625 40312
rect 367732 40205 367737 40312
rect 81365 39953 84874 40023
rect 84804 39583 84874 39953
rect 84801 39578 84874 39583
rect 84801 39518 84806 39578
rect 84866 39518 84874 39578
rect 84801 39513 84874 39518
rect 84804 39243 84874 39513
rect 84804 39238 84875 39243
rect 84804 39178 84810 39238
rect 84870 39178 84875 39238
rect 81027 39175 81093 39176
rect 80857 39171 81093 39175
rect 80857 39115 81032 39171
rect 81088 39115 81093 39171
rect 80857 39111 81093 39115
rect 81027 39110 81093 39111
rect 84804 39173 84875 39178
rect 84804 39031 84874 39173
rect 84801 39026 84874 39031
rect 84801 38966 84806 39026
rect 84866 38966 84874 39026
rect 84801 38961 84874 38966
rect 84804 38960 84874 38961
rect 80941 38578 81007 38581
rect 80839 38576 81012 38578
rect 80839 38520 80946 38576
rect 81002 38520 81012 38576
rect 80839 38518 81012 38520
rect 80941 38515 81007 38518
rect 16826 35740 32900 35880
rect 105589 35675 109435 35896
rect 244118 34975 246587 35026
rect 186561 34827 188561 34860
rect 10712 34600 20254 34726
rect 23902 34588 32518 34744
rect 134140 34561 134564 34696
rect 11216 34162 28318 34304
rect 186561 34181 186599 34827
rect 188523 34181 188561 34827
rect 192684 34699 193509 34834
rect 244118 34357 244169 34975
rect 246537 34357 246587 34975
rect 244118 34316 246587 34357
rect 186561 34153 188561 34181
rect 11700 33700 28318 33850
rect 229185 33665 231794 33754
rect 170217 33539 174718 33601
rect 12240 33310 20270 33474
rect 23930 33212 32120 33346
rect 229811 33305 231794 33394
rect 170873 33179 174718 33241
rect 15886 32884 31754 33018
rect 265730 32328 277810 32712
rect 280282 32380 284304 32764
rect 277072 32033 278516 32069
rect 232626 31763 234573 31847
rect 175028 31631 176381 31682
rect 175028 31064 175103 31631
rect 176317 31064 176381 31631
rect 232626 31208 232705 31763
rect 234494 31208 234573 31763
rect 277072 31714 277126 32033
rect 278462 31714 278516 32033
rect 277072 31675 278516 31714
rect 232626 31141 234573 31208
rect 175028 30976 176381 31064
rect 279429 30999 280873 31032
rect 279429 30680 279477 30999
rect 280813 30680 280873 30999
rect 279429 30638 280873 30680
rect 232626 29867 234573 29934
rect 175029 29713 176382 29766
rect 175029 29146 175090 29713
rect 176304 29146 176382 29713
rect 232626 29312 232722 29867
rect 234511 29312 234573 29867
rect 232626 29228 234573 29312
rect 175029 29060 176382 29146
rect 244359 29128 247187 29162
rect 186616 28962 188515 28995
rect 186616 28312 186663 28962
rect 188472 28312 188515 28962
rect 244359 28490 244399 29128
rect 247152 28490 247187 29128
rect 244359 28454 247187 28490
rect 186616 28284 188515 28312
rect 28884 28085 30639 28117
rect 28884 27838 29905 28085
rect 30580 27838 30639 28085
rect 28884 27797 30639 27838
rect 277097 26027 278517 26053
rect 257238 26004 257390 26022
rect 254078 25752 254748 25753
rect 257238 25752 257258 26004
rect 254078 25168 257258 25752
rect 12748 20078 20234 20232
rect 13270 19478 28314 19632
rect 13792 18878 24838 19032
rect 14268 18278 16804 18432
rect 105573 18024 109451 18261
rect 254078 17726 254748 25168
rect 257238 24982 257258 25168
rect 257372 24982 257390 26004
rect 277097 25773 277138 26027
rect 278478 25773 278517 26027
rect 277097 25742 278517 25773
rect 257238 24958 257390 24982
rect 279430 25119 280850 25144
rect 279430 24865 279469 25119
rect 280809 24865 280850 25119
rect 279430 24833 280850 24865
rect 255679 23915 257365 23995
rect 256050 23801 257365 23815
rect 256050 23745 257366 23801
rect 256050 23735 257365 23745
rect 265644 19318 277820 19702
rect 280320 19312 283544 19704
rect 367620 19696 367737 40205
rect 384352 39680 385786 39728
rect 384352 39126 384400 39680
rect 385734 39126 385786 39680
rect 384352 39078 385786 39126
rect 479068 38784 480580 41541
rect 479068 34694 479268 38784
rect 480424 34694 480580 38784
rect 479068 34472 480580 34694
rect 389683 32738 394881 32754
rect 389683 32467 389701 32738
rect 391045 32731 394881 32738
rect 391045 32474 393779 32731
rect 394848 32474 394881 32731
rect 391045 32467 394881 32474
rect 389683 32447 394881 32467
rect 430070 31895 433193 31918
rect 430070 31890 432505 31895
rect 430070 31573 430108 31890
rect 430715 31573 432505 31890
rect 430070 31571 432505 31573
rect 433161 31571 433193 31895
rect 430070 31545 433193 31571
rect 391405 29084 393015 29129
rect 391405 28593 391451 29084
rect 392975 28593 393015 29084
rect 391405 28550 393015 28593
rect 431742 22716 439077 22807
rect 431742 22602 432014 22716
rect 434717 22602 439077 22716
rect 431742 21785 431923 22602
rect 438850 21785 439077 22602
rect 472975 22662 478554 22814
rect 431742 21603 439077 21785
rect 464419 21999 464585 22012
rect 464419 21538 464430 21999
rect 464574 21538 464585 21999
rect 464419 21526 464585 21538
rect 464711 21998 464877 22012
rect 464711 21537 464722 21998
rect 464866 21537 464877 21998
rect 464711 21526 464877 21537
rect 465015 21997 465181 22012
rect 465015 21536 465027 21997
rect 465171 21536 465181 21997
rect 465015 21526 465181 21536
rect 465352 22001 465518 22013
rect 465352 21540 465360 22001
rect 465504 21540 465518 22001
rect 465352 21527 465518 21540
rect 467417 22000 467624 22011
rect 467417 21539 467428 22000
rect 467613 21539 467624 22000
rect 467417 21526 467624 21539
rect 472975 21637 473177 22662
rect 478353 21637 478554 22662
rect 472975 21503 478554 21637
rect 387791 21145 460622 21311
rect 430934 20715 459047 20886
rect 388429 20210 457482 20381
rect 388858 19819 455848 19990
rect 367620 19589 367625 19696
rect 367732 19589 367737 19696
rect 367620 19584 367737 19589
rect 386940 19448 451045 19619
rect 254078 17202 254104 17726
rect 254714 17202 254748 17726
rect 254078 17168 254748 17202
rect 294461 19081 295062 19197
rect 294461 16433 294545 19081
rect 295010 16433 295062 19081
rect 353180 18955 433270 19170
rect 436246 19036 446288 19220
rect 433055 18770 433270 18955
rect 386264 18510 430771 18718
rect 433055 18556 439885 18770
rect 433115 18555 439885 18556
rect 337270 17911 337370 18510
rect 417790 18122 417974 18370
rect 337270 17906 341158 17911
rect 337270 17816 341063 17906
rect 341153 17816 341158 17906
rect 337270 17811 341158 17816
rect 430563 17429 430771 18510
rect 439670 17463 439885 18555
rect 446062 17423 446288 19036
rect 450874 17354 451045 19448
rect 452474 18116 452676 19551
rect 454062 18112 454264 19028
rect 455677 17429 455848 19819
rect 457311 17411 457482 20210
rect 458876 17361 459047 20715
rect 460456 17376 460622 21145
rect 352777 17151 415493 17289
rect 353685 16561 415644 16728
rect 294461 16310 295062 16433
rect 4480 11266 4657 16241
rect 124105 12624 124487 12672
rect 90535 12520 90924 12560
rect 90535 10985 90573 12520
rect 90888 10985 90924 12520
rect 123574 11829 123957 11867
rect 90535 10924 90924 10985
rect 91072 11779 91458 11822
rect 91072 10993 91116 11779
rect 91423 10993 91458 11779
rect 91072 10933 91458 10993
rect 123574 10977 123624 11829
rect 123927 10977 123957 11829
rect 123574 10929 123957 10977
rect 124105 10975 124147 12624
rect 124449 10975 124487 12624
rect 124105 10928 124487 10975
rect 343299 9006 343429 14739
rect 343811 9306 343941 14739
rect 344323 9606 344453 14739
rect 344835 9906 344965 14739
rect 345347 10206 345477 14739
rect 345859 10506 345989 14739
rect 346371 10806 346501 14739
rect 346883 11106 347013 14739
rect 347395 11406 347525 14739
rect 348931 12306 349061 14739
rect 349443 12606 349573 14739
rect 349955 12906 350085 14739
rect 350467 13206 350597 14739
rect 350979 13506 351109 14739
rect 351491 13806 351621 14739
rect 351491 13666 354614 13806
rect 350979 13366 354078 13506
rect 350467 13066 353558 13206
rect 349955 12766 353048 12906
rect 349443 12466 352522 12606
rect 348931 12166 352018 12306
rect 347395 11266 350472 11406
rect 346883 10966 349940 11106
rect 346371 10666 349454 10806
rect 351878 10600 352018 12166
rect 352382 10702 352522 12466
rect 352908 10933 353048 12766
rect 353418 11285 353558 13066
rect 353938 11591 354078 13366
rect 354474 11859 354614 13666
rect 345859 10366 348916 10506
rect 345347 10066 348418 10206
rect 344835 9766 347898 9906
rect 344323 9466 347382 9606
rect 343811 9166 346868 9306
rect 343299 8866 346364 9006
rect 230142 8722 342687 8862
rect 13622 7878 252093 8006
rect 13622 7532 226852 7732
rect 345948 7494 354854 7890
rect 13622 7256 252093 7384
rect 13622 6910 226580 7110
rect 382141 7034 382261 7480
rect 468366 7245 468731 7264
rect 363174 7033 382261 7034
rect 363169 6931 382261 7033
rect 363174 6930 382261 6931
rect 468366 6914 468381 7245
rect 468715 7129 468731 7245
rect 482857 7129 482957 43639
rect 550355 35144 569352 35444
rect 527070 34320 535760 34532
rect 542818 34233 547933 34361
rect 548660 34195 555960 34323
rect 531337 33919 539216 34131
rect 548660 34011 548788 34195
rect 558400 34016 569956 34316
rect 542556 33883 548788 34011
rect 549285 33823 555613 33951
rect 549285 33702 549413 33823
rect 542024 33574 549413 33702
rect 528347 33278 535719 33506
rect 542299 33162 547651 33290
rect 550055 33232 570548 33532
rect 558128 27707 571158 28007
rect 526564 20541 535738 20719
rect 550056 20713 564520 21013
rect 558100 20100 565136 20400
rect 540888 17867 563742 18029
rect 540310 17502 563393 17664
rect 483374 8786 483515 14662
rect 483792 9224 483959 16171
rect 484194 9640 484333 17162
rect 538419 16757 565096 16884
rect 531374 16315 565746 16450
rect 530828 15869 566342 16022
rect 484527 10644 484647 15540
rect 487522 10794 488298 10844
rect 487522 10644 487572 10794
rect 484527 10524 487572 10644
rect 487522 10414 487572 10524
rect 488240 10414 488298 10794
rect 487522 10356 488298 10414
rect 484194 9501 555884 9640
rect 483792 9057 528101 9224
rect 555761 8952 555884 9501
rect 567984 9500 570458 9622
rect 555761 8829 562682 8952
rect 483374 8645 555532 8786
rect 555391 8441 555532 8645
rect 555391 8300 562143 8441
rect 563042 8429 571651 8552
rect 563545 8029 572311 8152
rect 492855 7629 564576 7752
rect 468715 7029 482957 7129
rect 468715 6914 468731 7029
rect 468366 6899 468731 6914
rect 13622 6635 555792 6762
rect 13622 6634 339282 6635
rect 340156 6634 555792 6635
rect 105723 6288 555792 6488
rect 105723 6012 555792 6140
rect 105723 5666 547764 5866
rect 105723 5390 547764 5518
rect 54 3500 20964 3538
rect 54 2550 20260 3500
rect 20922 2550 20964 3500
rect 54 2510 20964 2550
rect 557282 3138 572524 3168
rect 557282 2170 557330 3138
rect 557790 2170 572524 3138
rect 557282 2134 572524 2170
rect 21982 1143 256199 1291
rect 21982 843 256163 991
rect 22109 543 255792 691
rect 21982 243 256199 391
<< via3 >>
rect 508087 109535 508795 110004
rect 43650 106779 44525 107232
rect 509061 107636 509627 108138
rect 44952 105047 45825 105596
rect 90487 91240 90776 99164
rect 91536 91270 91825 99194
rect 96467 91204 96717 99138
rect 97389 91199 97639 99133
rect 120083 98530 121300 106035
rect 234448 104915 239019 106448
rect 118373 84581 120275 88705
rect 230496 84812 232362 85990
rect 28061 84214 30580 84482
rect 25531 83300 28093 83562
rect 142694 82140 143519 82275
rect 46174 80934 46578 81190
rect 159665 81202 160145 83248
rect 44940 80162 45820 80778
rect 141515 80655 142340 80790
rect 160460 80742 160761 82089
rect 160996 80732 161307 81841
rect 193329 81115 193632 81893
rect 193852 81115 194157 82259
rect 194429 81152 194994 83616
rect 207523 82259 208139 82413
rect 212513 80792 213299 80936
rect 46844 79704 47248 79960
rect 140440 79863 141141 80003
rect 198863 79994 199411 80135
rect 139559 79294 140240 79442
rect 203014 79434 203471 79576
rect 15440 78335 17907 78642
rect 43650 78584 44534 79042
rect 266396 91782 266692 94036
rect 267407 91782 267703 94036
rect 272379 91796 272620 94036
rect 273303 91819 273540 94027
rect 320963 91528 321227 93488
rect 321890 91560 322143 93472
rect 319004 88765 319323 90714
rect 319886 88736 320160 91499
rect 354382 101717 355624 106521
rect 465393 105291 467127 106993
rect 352789 84990 354530 91801
rect 498275 91530 498510 93854
rect 499190 91505 499425 93829
rect 504104 91513 504385 93849
rect 505121 91496 505402 93832
rect 554213 89107 555054 89337
rect 552725 88193 553869 88427
rect 473636 84830 475432 86252
rect 394019 80729 394553 83338
rect 394851 80687 395147 82606
rect 395370 80671 395671 81462
rect 427385 80611 427699 81409
rect 427915 80638 428234 82532
rect 428533 80656 429062 83660
rect 499949 82893 500235 84146
rect 501152 81984 501407 83150
rect 509068 82928 509620 83514
rect 545974 82338 546865 83115
rect 508114 81348 508775 82112
rect 450757 80161 451373 80303
rect 375497 79999 376097 80126
rect 374700 79434 375223 79563
rect 451681 79499 452277 79631
rect 543189 79844 544669 80189
rect 566647 83208 567525 83547
rect 562875 82178 563960 82526
rect 20283 77294 22755 77609
rect 7360 64720 8556 65236
rect 11043 64365 14614 65195
rect 132948 60752 133712 61258
rect 414932 60678 415612 61829
rect 153572 59658 155089 60010
rect 29923 56030 30568 56270
rect 25084 55113 25761 55346
rect 130264 58260 130786 59100
rect 150103 59034 151655 59383
rect 183998 59273 185192 59797
rect 212513 59792 214046 60138
rect 209089 59178 210622 59524
rect 405465 59616 406501 59916
rect 189798 58319 190768 58513
rect 129052 57232 129570 58028
rect 130252 56262 130774 56982
rect 131492 55114 132264 56024
rect 342211 55198 342363 56112
rect 342515 55217 342664 56109
rect 352180 58638 353960 59225
rect 372341 58463 373424 59420
rect 529578 57678 529863 58947
rect 530611 57726 530896 58995
rect 535562 58682 535808 59924
rect 536487 58686 536733 59928
rect 132702 54136 133477 54865
rect 191120 54832 192099 55017
rect 132724 52870 133492 53942
rect 182438 52513 183994 52696
rect 186566 52384 187774 52604
rect 374345 52579 375302 52920
rect 421070 51773 421767 51919
rect 15441 50156 16081 50456
rect 131501 49554 132272 50210
rect 20278 49121 20906 49409
rect 86040 48708 86615 49374
rect 364765 49357 364915 50211
rect 368319 49227 369200 49395
rect 421046 48341 421743 48487
rect 130254 46352 130776 47192
rect 420803 47023 421743 47148
rect 129052 45292 129564 46104
rect 420789 46034 421670 46173
rect 130246 44332 130791 45079
rect 402922 44613 403374 45342
rect 403806 44919 404042 45940
rect 81394 43170 82156 44114
rect 29917 42025 30568 42289
rect 99918 42201 100644 42962
rect 25082 41122 25759 41355
rect 82822 40922 83516 41778
rect 562759 60236 564261 60665
rect 566623 58523 567534 59030
rect 551991 54794 552467 55050
rect 553227 53876 553703 54132
rect 556070 48910 556495 49239
rect 557345 47868 557770 48197
rect 385274 43242 386087 43716
rect 452319 41819 459350 42872
rect 384078 41169 385891 41614
rect 15443 36154 16083 36454
rect 20279 35128 20907 35416
rect 186599 34181 188523 34827
rect 244169 34357 246537 34975
rect 175103 31064 176317 31631
rect 232705 31208 234494 31763
rect 277126 31714 278462 32033
rect 279477 30680 280813 30999
rect 175090 29146 176304 29713
rect 232722 29312 232969 29867
rect 232969 29312 234511 29867
rect 186663 28312 188472 28962
rect 244399 28490 247152 29128
rect 29905 27838 30580 28085
rect 25087 26929 25764 27162
rect 15423 21969 16096 22246
rect 20266 20930 20894 21218
rect 277138 25773 278478 26027
rect 279469 24865 280809 25119
rect 384400 39126 385734 39680
rect 479268 34694 480424 38784
rect 389701 32467 391045 32738
rect 432505 31571 433161 31895
rect 391451 28615 392065 29084
rect 392065 28615 392969 29084
rect 392969 28615 392975 29084
rect 391451 28593 392975 28615
rect 432014 22602 434717 22716
rect 432014 21830 434717 22602
rect 473177 21637 478353 22662
rect 254104 17202 254714 17726
rect 294545 16433 295010 19081
rect 341612 14571 341779 15785
rect 341910 14571 342077 15785
rect 90573 10985 90888 12520
rect 91116 10993 91423 11779
rect 123624 10977 123927 11829
rect 124147 10975 124449 12624
rect 148560 9670 149640 10004
rect 207488 9803 208597 10148
rect 156146 9104 157226 9438
rect 215049 9233 216158 9578
rect 457704 6898 458043 7228
rect 468381 6914 468715 7245
rect 533708 41736 534074 41995
rect 552005 41575 552430 41808
rect 532870 40806 533236 41065
rect 553252 40643 553677 40876
rect 537333 35840 537724 36166
rect 556063 35680 556515 35981
rect 536094 34797 536485 35123
rect 557338 34631 557790 34932
rect 533717 28161 534113 28437
rect 551998 28194 552437 28406
rect 532860 27232 533256 27508
rect 553259 27275 553698 27515
rect 537335 22277 537727 22596
rect 556049 22285 556515 22600
rect 536097 21250 536489 21569
rect 557324 21277 557790 21592
rect 487572 10414 488240 10794
rect 20260 2550 20922 3500
rect 557330 2170 557790 3138
<< metal4 >>
rect 8212 112722 8412 115349
rect 8812 113266 9012 115200
rect 32212 112726 32412 115349
rect 32812 113720 33012 115200
rect 56212 112718 56412 115349
rect 56812 114060 57012 115200
rect 80212 112730 80412 115349
rect 80812 114400 81012 115200
rect 115352 113486 120228 115192
rect 93932 112283 120228 113486
rect 120452 112283 125328 115192
rect 150212 112722 150412 115349
rect 150812 113004 151012 115200
rect 174212 112790 174412 115349
rect 174812 113454 175012 115200
rect 198212 112730 198412 115349
rect 198812 113850 199012 115200
rect 222212 112722 222412 115349
rect 222812 114216 223012 115200
rect 43628 107232 44554 107283
rect 43628 106779 43650 107232
rect 44525 106779 44554 107232
rect 5430 90172 5580 92568
rect 5430 71238 5580 89609
rect 4544 16040 4669 63491
rect 6068 50265 6218 76949
rect 6568 29220 6718 76520
rect 7711 68897 7989 93595
rect 15396 78676 16135 91034
rect 15393 78642 17975 78676
rect 15393 78335 15440 78642
rect 17907 78335 17975 78642
rect 15393 78297 17975 78335
rect 15396 74356 16135 78297
rect 20222 77664 20961 91034
rect 25048 84356 25787 91034
rect 29874 84506 30613 91034
rect 25048 82430 25090 84356
rect 25749 83592 25787 84356
rect 28033 84482 30615 84506
rect 28033 84214 28061 84482
rect 30580 84214 30615 84482
rect 28033 84191 30615 84214
rect 25749 83562 28129 83592
rect 28093 83300 28129 83562
rect 25749 83270 28129 83300
rect 25749 82430 25787 83270
rect 20220 77609 22806 77664
rect 20220 77294 20283 77609
rect 22755 77294 22806 77609
rect 20220 77264 22806 77294
rect 15396 69442 15421 74356
rect 16093 69442 16135 74356
rect 7293 65236 8639 68897
rect 7293 64720 7360 65236
rect 8556 64720 8639 65236
rect 7293 64686 8639 64720
rect 6956 64408 8639 64686
rect 10917 65195 14755 65344
rect 6956 30236 7234 64408
rect 10917 64365 11043 65195
rect 14614 64365 14755 65195
rect 10917 64208 14755 64365
rect 7636 15548 7764 61890
rect 368 15420 7764 15548
rect 108 0 236 3538
rect 368 0 496 15420
rect 8148 15036 8276 61506
rect 15396 50456 16135 69442
rect 15396 50156 15441 50456
rect 16081 50156 16135 50456
rect 880 14908 8276 15036
rect 620 0 748 3538
rect 880 0 1008 14908
rect 8660 14524 8788 48786
rect 1392 14396 8788 14524
rect 1132 0 1260 3538
rect 1392 0 1520 14396
rect 9172 14012 9300 48340
rect 1904 13884 9300 14012
rect 1644 0 1772 3538
rect 1904 0 2032 13884
rect 9684 13500 9812 47862
rect 2416 13372 9812 13500
rect 2156 0 2284 3538
rect 2416 0 2544 13372
rect 10196 12988 10324 47496
rect 15396 36454 16135 50156
rect 15396 36154 15443 36454
rect 16083 36154 16135 36454
rect 2928 12860 10324 12988
rect 2668 0 2796 3538
rect 2928 0 3056 12860
rect 10708 12476 10836 34772
rect 3440 12348 10836 12476
rect 3180 0 3308 3538
rect 3440 0 3568 12348
rect 11220 11964 11348 34318
rect 3952 11836 11348 11964
rect 3692 0 3820 3538
rect 3952 0 4080 11836
rect 4204 0 4332 3538
rect 4464 0 4592 11398
rect 11744 10940 11872 33880
rect 4976 10812 11872 10940
rect 4716 0 4844 3538
rect 4976 0 5104 10812
rect 12256 10428 12384 33494
rect 15396 22246 16135 36154
rect 15396 21969 15423 22246
rect 16096 21969 16135 22246
rect 15396 20749 16135 21969
rect 20222 67331 20961 77264
rect 20222 62506 20258 67331
rect 20918 62506 20961 67331
rect 20222 49409 20961 62506
rect 20222 49121 20278 49409
rect 20906 49121 20961 49409
rect 20222 35416 20961 49121
rect 20222 35128 20279 35416
rect 20907 35128 20961 35416
rect 20222 21218 20961 35128
rect 20222 20930 20266 21218
rect 20894 20930 20961 21218
rect 5488 10300 12384 10428
rect 5228 0 5356 3538
rect 5488 0 5616 10300
rect 12768 9916 12896 20320
rect 6000 9788 12896 9916
rect 5740 0 5868 3538
rect 6000 0 6128 9788
rect 13280 9404 13408 19680
rect 6512 9276 13408 9404
rect 6252 0 6380 3538
rect 6512 0 6640 9276
rect 13780 7048 13908 19112
rect 14280 7696 14408 18452
rect 6772 0 6900 3538
rect 20222 3500 20961 20930
rect 25048 55346 25787 82430
rect 25048 55113 25084 55346
rect 25761 55113 25787 55346
rect 25048 41355 25787 55113
rect 25048 41122 25082 41355
rect 25759 41122 25787 41355
rect 25048 27162 25787 41122
rect 25048 26929 25087 27162
rect 25764 26929 25787 27162
rect 25048 20839 25787 26929
rect 29874 80360 30613 84191
rect 29874 78434 29921 80360
rect 30580 78434 30613 80360
rect 29874 56270 30613 78434
rect 31520 72112 31660 76956
rect 31920 72596 32060 78092
rect 32320 73104 32460 89140
rect 32720 73612 32860 89562
rect 34700 77190 35439 90407
rect 37765 84315 38436 84405
rect 37765 82462 37821 84315
rect 38379 82462 38436 84315
rect 37765 82407 38436 82462
rect 34700 76451 37696 77190
rect 36957 74322 37696 76451
rect 29874 56030 29923 56270
rect 30568 56030 30613 56270
rect 29874 42289 30613 56030
rect 29874 42025 29917 42289
rect 30568 42025 30613 42289
rect 29874 28085 30613 42025
rect 31540 32164 31680 66050
rect 31940 33284 32080 66558
rect 32340 34580 32480 67064
rect 32740 35722 32880 67600
rect 33140 46976 33280 68100
rect 33540 47218 33680 68614
rect 33940 48620 34080 70178
rect 34340 49708 34480 70650
rect 34736 60564 34876 71166
rect 35140 61122 35280 71638
rect 36957 69435 37010 74322
rect 37641 69435 37696 74322
rect 36957 69381 37696 69435
rect 38031 60763 38428 82407
rect 38635 80323 39312 80391
rect 38635 78461 38721 80323
rect 39238 78461 39312 80323
rect 38635 78385 39312 78461
rect 36019 60366 38428 60763
rect 36019 56651 36416 60366
rect 38764 60041 39141 78385
rect 39526 67339 40265 91073
rect 43628 79042 44554 106779
rect 43628 78584 43650 79042
rect 44534 78584 44554 79042
rect 40715 74380 41327 74393
rect 39526 62500 39559 67339
rect 40217 62500 40265 67339
rect 39526 62440 40265 62500
rect 40704 74319 41327 74380
rect 40704 69472 40801 74319
rect 41224 69472 41327 74319
rect 40704 69394 41327 69472
rect 43628 74274 44554 78584
rect 43628 69482 43708 74274
rect 44464 69482 44554 74274
rect 36493 59664 39141 60041
rect 36493 56651 36870 59664
rect 40704 59512 41078 69394
rect 43628 69340 44554 69482
rect 44922 105596 45848 105668
rect 44922 105047 44952 105596
rect 45825 105047 45848 105596
rect 44922 80778 45848 105047
rect 91063 104437 91223 106450
rect 89948 104277 91228 104437
rect 46720 84312 47326 84388
rect 46720 82470 46784 84312
rect 47234 82470 47326 84312
rect 46720 82394 47326 82470
rect 44922 80162 44940 80778
rect 45820 80162 45848 80778
rect 46160 81190 46604 81232
rect 46160 80934 46174 81190
rect 46578 80934 46604 81190
rect 46160 80888 46604 80934
rect 46160 80480 46608 80888
rect 41453 67339 42060 67417
rect 41453 62466 41507 67339
rect 42011 62466 42060 67339
rect 41453 62396 42060 62466
rect 44922 67310 45848 80162
rect 46094 80306 46700 80480
rect 46094 78464 46174 80306
rect 46624 78464 46700 80306
rect 46830 79960 47274 82394
rect 46830 79704 46844 79960
rect 47248 79704 47274 79960
rect 46830 79658 47274 79704
rect 46094 78394 46700 78464
rect 89534 76256 89694 98060
rect 89948 76700 90108 104277
rect 90411 99164 90852 99255
rect 90411 91240 90487 99164
rect 90776 91240 90852 99164
rect 90411 81704 90852 91240
rect 91460 99194 91901 99240
rect 91460 91270 91536 99194
rect 91825 91270 91901 99194
rect 91460 82749 91901 91270
rect 91460 82308 92344 82749
rect 90411 81263 91354 81704
rect 44922 62518 45004 67310
rect 45760 62518 45848 67310
rect 64372 63460 65022 74480
rect 74350 70632 74519 74403
rect 83820 74312 84682 74510
rect 83820 69498 83914 74312
rect 84573 69498 84682 74312
rect 85180 70078 85349 74403
rect 44922 62414 45848 62518
rect 36952 59138 41078 59512
rect 36952 56583 37326 59138
rect 41457 58874 41818 62396
rect 37441 58513 41818 58874
rect 83820 61116 84682 69498
rect 90913 67357 91354 81263
rect 91903 74308 92344 82308
rect 91903 69425 91979 74308
rect 92280 69425 92344 74308
rect 91903 69372 92344 69425
rect 83820 58740 83875 61116
rect 84621 58740 84682 61116
rect 37441 56583 37802 58513
rect 81366 44114 82186 46112
rect 81366 43170 81394 44114
rect 82156 43170 82186 44114
rect 29874 27838 29905 28085
rect 30580 27838 30613 28085
rect 29874 21025 30613 27838
rect 81366 13352 82186 43170
rect 82794 41778 83552 41845
rect 82794 40922 82822 41778
rect 83516 40922 83552 41778
rect 81366 13322 82376 13352
rect 81254 13072 82376 13322
rect 81254 11629 81321 13072
rect 82276 11629 82376 13072
rect 81254 11567 82376 11629
rect 82794 9768 83552 40922
rect 83820 36986 84682 58740
rect 85014 67220 85891 67329
rect 85014 62454 85099 67220
rect 85769 62454 85891 67220
rect 85014 38291 85891 62454
rect 90913 62474 90989 67357
rect 91290 62474 91354 67357
rect 90913 62409 91354 62474
rect 93932 49454 94704 112283
rect 99902 111535 99996 111536
rect 120452 111535 122738 112283
rect 99902 110414 122738 111535
rect 131293 111807 132395 111935
rect 96373 99138 96814 99240
rect 96373 91204 96467 99138
rect 96717 91204 96814 99138
rect 96373 84319 96814 91204
rect 96373 82461 96440 84319
rect 96740 82461 96814 84319
rect 96373 82386 96814 82461
rect 97286 99133 97727 99255
rect 97286 91199 97389 99133
rect 97639 91199 97727 99133
rect 97286 80304 97727 91199
rect 97286 78446 97352 80304
rect 97652 78446 97727 80304
rect 97286 78359 97727 78446
rect 85977 49374 94704 49454
rect 85977 48708 86040 49374
rect 86615 48708 94704 49374
rect 85977 48682 94704 48708
rect 99902 42962 100674 110414
rect 131293 110345 131380 111807
rect 132311 110345 132395 111807
rect 131293 110136 132395 110345
rect 102886 77106 103046 106204
rect 119630 106035 121653 106475
rect 119630 98530 120083 106035
rect 121300 98530 121653 106035
rect 103924 77486 104084 98184
rect 119630 94542 121653 98530
rect 119630 92519 123743 94542
rect 118187 88705 120438 88927
rect 118187 84581 118373 88705
rect 120275 84581 120438 88705
rect 118187 74180 120438 84581
rect 118187 69535 118373 74180
rect 120308 69535 120438 74180
rect 118187 69368 120438 69535
rect 121720 67196 123743 92519
rect 130216 84334 130820 84412
rect 130216 82434 130258 84334
rect 130778 82434 130820 84334
rect 129008 80342 129612 80448
rect 129008 78442 129052 80342
rect 129572 78442 129612 80342
rect 127660 74293 128447 74395
rect 127660 69488 127814 74293
rect 128339 69488 128447 74293
rect 121720 62593 121918 67196
rect 123526 62593 123743 67196
rect 121720 62313 123743 62593
rect 126351 67298 127121 67453
rect 126351 62493 126488 67298
rect 127013 62493 127121 67298
rect 99902 42201 99918 42962
rect 100644 42201 100674 42962
rect 99902 42079 100674 42201
rect 85014 37414 89915 38291
rect 126351 38053 127121 62493
rect 83820 36124 89059 36986
rect 89492 36490 89915 37414
rect 125096 37372 127121 38053
rect 125096 36600 125525 37372
rect 127660 36945 128447 69488
rect 129008 58028 129612 78442
rect 129008 57232 129052 58028
rect 129570 57232 129612 58028
rect 129008 46104 129612 57232
rect 129008 45292 129052 46104
rect 129564 45292 129612 46104
rect 129008 45150 129612 45292
rect 130216 59100 130820 82434
rect 130216 58260 130264 59100
rect 130786 58260 130820 59100
rect 130216 56982 130820 58260
rect 130216 56262 130252 56982
rect 130774 56262 130820 56982
rect 131552 57218 132395 110136
rect 132904 109413 134006 109537
rect 132904 107951 132983 109413
rect 133914 107951 134006 109413
rect 132904 107734 134006 107951
rect 132904 61258 133750 107734
rect 234318 106448 239118 115200
rect 244018 111534 248818 115200
rect 258277 111534 259374 112898
rect 265212 112718 265412 115349
rect 265812 114806 266012 115200
rect 244018 106734 262452 111534
rect 234318 104915 234448 106448
rect 239019 104915 239118 106448
rect 139541 84335 140260 84392
rect 139541 82437 139578 84335
rect 140216 82437 140260 84335
rect 139541 79442 140260 82437
rect 142675 82275 143534 82316
rect 142675 82140 142694 82275
rect 143519 82140 143534 82275
rect 141495 80790 142375 80857
rect 141495 80655 141515 80790
rect 142340 80655 142375 80790
rect 139541 79294 139559 79442
rect 140240 79294 140260 79442
rect 139541 79272 140260 79294
rect 140423 80339 141167 80392
rect 140423 80003 140461 80339
rect 141130 80003 141167 80339
rect 140423 79863 140440 80003
rect 141141 79863 141167 80003
rect 140423 78428 140461 79863
rect 141130 78428 141167 79863
rect 140423 78389 141167 78428
rect 141495 74335 142375 80655
rect 141495 69463 141534 74335
rect 142314 69463 142375 74335
rect 141495 69351 142375 69463
rect 142675 67337 143534 82140
rect 154799 80342 155260 90399
rect 155587 84353 156070 88858
rect 155587 82449 155647 84353
rect 156028 82449 156070 84353
rect 155587 82412 156070 82449
rect 154799 78438 154843 80342
rect 155224 78438 155260 80342
rect 154799 78396 155260 78438
rect 156483 76251 156623 92461
rect 155743 76111 156623 76251
rect 153550 74319 155115 74426
rect 153550 69472 153620 74319
rect 155025 69472 155115 74319
rect 142675 62453 142726 67337
rect 143472 62453 143534 67337
rect 142675 62396 143534 62453
rect 150076 67300 151681 67393
rect 150076 62514 150178 67300
rect 151580 62514 151681 67300
rect 132904 60752 132948 61258
rect 133712 60752 133750 61258
rect 132904 60662 133750 60752
rect 150076 59383 151681 62514
rect 153550 60010 155115 69472
rect 155743 62443 155883 76111
rect 157083 71615 157223 93935
rect 157683 71054 157823 95236
rect 160964 84342 161341 84383
rect 159562 83248 160245 83335
rect 158598 76445 159218 81229
rect 159562 81202 159665 83248
rect 160145 81202 160245 83248
rect 160964 82456 161026 84342
rect 161275 82456 161341 84342
rect 160429 82141 160805 82143
rect 159562 77834 160245 81202
rect 160428 82089 160805 82141
rect 160428 80742 160460 82089
rect 160761 80742 160805 82089
rect 160964 81881 161341 82456
rect 160428 80685 160805 80742
rect 160959 81841 161341 81881
rect 160959 80732 160996 81841
rect 161307 80732 161341 81841
rect 160959 80688 161341 80732
rect 160428 80335 160804 80685
rect 160964 80683 161341 80688
rect 182457 84328 183291 84416
rect 182457 82473 182529 84328
rect 183204 82473 183291 84328
rect 160428 78449 160495 80335
rect 160744 78449 160804 80335
rect 160428 78395 160804 78449
rect 159562 77151 160754 77834
rect 158598 75586 159834 76445
rect 159214 74294 159834 75586
rect 159214 69523 159333 74294
rect 159746 69523 159834 74294
rect 159214 69406 159834 69523
rect 160071 67284 160754 77151
rect 160071 62500 160173 67284
rect 160653 62500 160754 67284
rect 160071 62386 160754 62500
rect 153550 59658 153572 60010
rect 155089 59658 155115 60010
rect 153550 59623 155115 59658
rect 150076 59034 150103 59383
rect 151655 59034 151681 59383
rect 150076 58995 151681 59034
rect 131552 56375 133516 57218
rect 130216 47192 130820 56262
rect 130216 46352 130254 47192
rect 130776 46352 130820 47192
rect 130216 45079 130820 46352
rect 130216 44332 130246 45079
rect 130791 44332 130820 45079
rect 130216 44285 130820 44332
rect 131454 56024 132316 56114
rect 131454 55114 131492 56024
rect 132264 55114 132316 56024
rect 131454 50210 132316 55114
rect 132673 54865 133516 56375
rect 132673 54136 132702 54865
rect 133477 54136 133516 54865
rect 132673 54101 133516 54136
rect 131454 49554 131501 50210
rect 132272 49554 132316 50210
rect 125663 36158 128447 36945
rect 82680 9706 83552 9768
rect 90535 12520 90924 12560
rect 90535 10985 90573 12520
rect 90888 10985 90924 12520
rect 82680 9464 83802 9706
rect 82680 8021 82751 9464
rect 83706 8021 83802 9464
rect 82680 7933 83802 8021
rect 20222 2550 20260 3500
rect 20922 2550 20961 3500
rect 20222 2509 20961 2550
rect 90535 2234 90924 10985
rect 91072 11779 91458 11822
rect 91072 10993 91116 11779
rect 91423 10993 91458 11779
rect 91072 10933 91458 10993
rect 91072 4643 91454 10933
rect 106490 6470 106773 18150
rect 108128 5864 108411 35848
rect 124105 12624 124487 12672
rect 123574 11829 123957 11867
rect 123574 10977 123624 11829
rect 123927 10977 123957 11829
rect 91072 3174 91118 4643
rect 91406 3174 91454 4643
rect 91072 3123 91454 3174
rect 123574 4661 123957 10977
rect 123574 3181 123625 4661
rect 123912 3181 123957 4661
rect 123574 3128 123957 3181
rect 124105 10975 124147 12624
rect 124449 10975 124487 12624
rect 90535 765 90590 2234
rect 90878 765 90924 2234
rect 90535 694 90924 765
rect 124105 2237 124487 10975
rect 131454 7246 132316 49554
rect 132676 53942 133538 53999
rect 132676 52870 132724 53942
rect 133492 52870 133538 53942
rect 132676 9650 133538 52870
rect 182457 52741 183291 82473
rect 193282 84330 193664 84390
rect 193282 82436 193333 84330
rect 193619 82436 193664 84330
rect 193282 81893 193664 82436
rect 194372 83616 195054 83685
rect 193282 81115 193329 81893
rect 193632 81115 193664 81893
rect 193282 81070 193664 81115
rect 193813 82259 194192 82310
rect 193813 81115 193852 82259
rect 194157 81115 194192 82259
rect 184069 80307 185166 80411
rect 184069 78472 184167 80307
rect 185074 78472 185166 80307
rect 184069 59846 185166 78472
rect 186678 80328 187330 80423
rect 186678 78451 186750 80328
rect 187269 78451 187330 80328
rect 183932 59797 185250 59846
rect 183932 59273 183998 59797
rect 185192 59273 185250 59797
rect 183932 59224 185250 59273
rect 182377 52696 184035 52741
rect 182377 52513 182438 52696
rect 183994 52513 184035 52696
rect 186678 52655 187330 78451
rect 193813 80343 194192 81115
rect 193813 78449 193869 80343
rect 194155 78449 194192 80343
rect 193813 78388 194192 78449
rect 194372 81152 194429 83616
rect 194994 81152 195054 83616
rect 191197 74303 191960 74435
rect 191197 69495 191297 74303
rect 191872 69495 191960 74303
rect 189900 67303 190646 67404
rect 189900 62495 189982 67303
rect 190557 62495 190646 67303
rect 189900 58535 190646 62495
rect 189741 58513 190803 58535
rect 189741 58319 189798 58513
rect 190768 58319 190803 58513
rect 189741 58275 190803 58319
rect 182377 52464 184035 52513
rect 186469 52604 187820 52655
rect 186469 52451 186566 52604
rect 186479 52384 186566 52451
rect 187774 52384 187820 52604
rect 186479 52333 187820 52384
rect 189900 34970 190646 58275
rect 191197 55048 191960 69495
rect 194372 67249 195054 81152
rect 195402 74320 196022 81692
rect 195402 69507 195491 74320
rect 195955 69507 196022 74320
rect 197189 72129 197329 95496
rect 197789 72665 197929 94195
rect 198389 76286 198529 92721
rect 198846 80358 199427 90554
rect 199813 84345 200411 89132
rect 230333 85990 232507 86189
rect 230333 84812 230496 85990
rect 232362 84812 232507 85990
rect 199813 82511 199850 84345
rect 200371 82511 200411 84345
rect 199813 82451 200411 82511
rect 202995 84336 203490 84397
rect 198846 80135 198882 80358
rect 199386 80135 199427 80358
rect 198846 79994 198863 80135
rect 199411 79994 199427 80135
rect 198846 78457 198882 79994
rect 199386 78457 199427 79994
rect 202995 82447 203025 84336
rect 203443 82447 203490 84336
rect 202995 79576 203490 82447
rect 202995 79434 203014 79576
rect 203471 79434 203490 79576
rect 202995 79420 203490 79434
rect 207511 82413 208154 82430
rect 207511 82259 207523 82413
rect 208139 82259 208154 82413
rect 198846 78407 199427 78457
rect 198389 76146 199643 76286
rect 195402 69404 196022 69507
rect 194372 62511 194459 67249
rect 194939 62511 195054 67249
rect 199503 62798 199643 76146
rect 207511 67295 208154 82259
rect 212491 80936 213326 80968
rect 212491 80792 212513 80936
rect 213299 80792 213326 80936
rect 212491 74394 213326 80792
rect 212482 74261 214090 74394
rect 212482 69514 212614 74261
rect 213958 69514 214090 74261
rect 194372 62393 195054 62511
rect 207511 62469 207583 67295
rect 208056 62469 208154 67295
rect 207511 62401 208154 62469
rect 209061 67252 210661 67393
rect 209061 62505 209202 67252
rect 210546 62505 210661 67252
rect 209061 59524 210661 62505
rect 212482 60138 214090 69514
rect 228882 67552 229022 78168
rect 230333 74231 232507 84812
rect 230333 69592 230551 74231
rect 232344 69592 232507 74231
rect 230333 69501 232507 69592
rect 230333 69339 232508 69501
rect 231782 69338 232508 69339
rect 228882 67412 230126 67552
rect 212482 59792 212513 60138
rect 214046 59792 214090 60138
rect 212482 59764 214090 59792
rect 209061 59178 209089 59524
rect 210622 59178 210661 59524
rect 209061 59110 210661 59178
rect 191072 55017 192134 55048
rect 191072 54832 191120 55017
rect 192099 54832 192134 55017
rect 191072 54788 192134 54832
rect 186484 34827 190646 34970
rect 186484 34224 186599 34827
rect 186561 34181 186599 34224
rect 188523 34224 190646 34827
rect 188523 34181 188561 34224
rect 186561 34153 188561 34181
rect 172180 31631 176391 31718
rect 172180 31064 175103 31631
rect 176317 31064 176391 31631
rect 172180 30956 176391 31064
rect 132676 8142 132718 9650
rect 133480 8142 133538 9650
rect 132676 8083 133538 8142
rect 137668 7520 137905 10979
rect 131454 5738 131510 7246
rect 132272 5738 132316 7246
rect 138033 6919 138270 10571
rect 148524 10004 149674 10045
rect 148524 9670 148560 10004
rect 149640 9670 149674 10004
rect 131454 5674 132316 5738
rect 124105 757 124153 2237
rect 124440 757 124487 2237
rect 124105 709 124487 757
rect 148524 2183 149674 9670
rect 156106 9438 157265 9512
rect 156106 9104 156146 9438
rect 157226 9104 157265 9438
rect 156106 4622 157265 9104
rect 166832 6960 167058 10596
rect 167200 7625 167426 11017
rect 156106 3258 156181 4622
rect 157163 3258 157265 4622
rect 156106 3137 157265 3258
rect 148524 819 148608 2183
rect 149590 819 149674 2183
rect 148524 716 149674 819
rect 172180 2245 172942 30956
rect 172180 759 172217 2245
rect 172892 759 172942 2245
rect 172180 582 172942 759
rect 173380 29713 176454 29784
rect 173380 29146 175090 29713
rect 176304 29146 176454 29713
rect 173380 29022 176454 29146
rect 191197 29022 191960 54788
rect 173380 4662 174142 29022
rect 186561 28962 191960 29022
rect 186561 28312 186663 28962
rect 188472 28312 191960 28962
rect 186561 28259 191960 28312
rect 196636 7541 196852 10645
rect 196990 7035 197206 10636
rect 207459 10148 208632 10201
rect 207459 9803 207488 10148
rect 208597 9803 208632 10148
rect 173380 3176 173431 4662
rect 174106 3176 174142 4662
rect 173380 582 174142 3176
rect 207459 2191 208632 9803
rect 215017 9578 216181 9670
rect 215017 9233 215049 9578
rect 216158 9233 216181 9578
rect 215017 4611 216181 9233
rect 225800 6956 226016 10641
rect 226149 7562 226365 10828
rect 229986 8741 230126 67412
rect 234318 67234 239118 104915
rect 247351 74305 248551 74488
rect 247351 69468 247420 74305
rect 248462 69468 248551 74305
rect 234318 62540 234444 67234
rect 238960 62540 239118 67234
rect 234318 62260 239118 62540
rect 245387 67297 246556 67450
rect 245387 62489 245474 67297
rect 246432 62489 246556 67297
rect 245387 35277 246556 62489
rect 244055 35026 246556 35277
rect 244055 34975 246587 35026
rect 244055 34357 244169 34975
rect 246537 34357 246587 34975
rect 244055 34316 246587 34357
rect 244055 34108 246556 34316
rect 230480 31763 234623 31876
rect 230480 31208 232705 31763
rect 234494 31208 234623 31763
rect 230480 31114 234623 31208
rect 215017 3227 215109 4611
rect 216072 3227 216181 4611
rect 215017 3126 216181 3227
rect 207459 807 207569 2191
rect 208532 807 208632 2191
rect 207459 697 208632 807
rect 230480 2250 231242 31114
rect 230480 759 230517 2250
rect 231189 759 231242 2250
rect 230480 582 231242 759
rect 231680 29867 234634 29973
rect 231680 29312 232722 29867
rect 234511 29312 234634 29867
rect 247351 29441 248551 69468
rect 253253 74267 256464 74389
rect 253253 69491 253359 74267
rect 256333 69491 256464 74267
rect 231680 29211 234634 29312
rect 231680 4664 232442 29211
rect 244288 29128 248551 29441
rect 244288 28490 244399 29128
rect 247152 28490 248551 29128
rect 244288 28241 248551 28490
rect 249302 67270 252513 67473
rect 249302 62494 249437 67270
rect 252411 62494 252513 67270
rect 249302 22684 252513 62494
rect 253253 38560 256464 69491
rect 257299 74319 257781 74472
rect 257299 69460 257364 74319
rect 257711 69460 257781 74319
rect 257299 61653 257781 69460
rect 258452 67274 262452 106734
rect 266333 94036 266733 94082
rect 266333 91782 266396 94036
rect 266692 91782 266733 94036
rect 266333 79638 266733 91782
rect 267362 94036 267762 94082
rect 267362 91782 267407 94036
rect 267703 91782 267762 94036
rect 267362 81062 267762 91782
rect 272334 94036 272652 94073
rect 272334 91796 272379 94036
rect 272620 91796 272652 94036
rect 268455 84351 268937 84489
rect 268455 82442 268502 84351
rect 268889 82442 268937 84351
rect 267362 80662 268037 81062
rect 266333 79238 267198 79638
rect 258452 62522 258542 67274
rect 262334 62522 262452 67274
rect 258452 62260 262452 62522
rect 257299 61171 259916 61653
rect 263920 61115 264402 67375
rect 266798 67328 267198 79238
rect 267637 74348 268037 80662
rect 267637 69489 267689 74348
rect 267990 69489 268037 74348
rect 267637 69416 268037 69489
rect 266798 62501 266840 67328
rect 267165 62501 267198 67328
rect 266798 62443 267198 62501
rect 268455 61155 268937 82442
rect 272334 84387 272652 91796
rect 273262 94027 273580 94069
rect 273262 91819 273303 94027
rect 273540 91819 273580 94027
rect 272334 84347 272678 84387
rect 272334 82464 272385 84347
rect 272639 82464 272678 84347
rect 272334 82400 272678 82464
rect 272336 82386 272678 82400
rect 273262 80533 273580 91819
rect 272983 80334 273580 80533
rect 272983 78456 273026 80334
rect 273529 78456 273580 80334
rect 272983 78403 273580 78456
rect 272983 60890 273465 78403
rect 277487 74336 277969 74510
rect 277487 69450 277546 74336
rect 277912 69450 277969 74336
rect 275075 67273 275798 67409
rect 275075 62522 275169 67273
rect 275693 62522 275798 67273
rect 275075 41647 275798 62522
rect 277487 60874 277969 69450
rect 279782 74306 280505 74464
rect 279782 69470 279860 74306
rect 280452 69470 280505 74306
rect 275075 40924 278059 41647
rect 253253 35349 257654 38560
rect 277336 32069 278059 40924
rect 277072 32033 278516 32069
rect 277072 31714 277126 32033
rect 278462 31714 278516 32033
rect 277072 31675 278516 31714
rect 279782 31032 280505 69470
rect 282035 67330 282517 67464
rect 282035 62444 282083 67330
rect 282449 62444 282517 67330
rect 282035 60929 282517 62444
rect 279429 30999 280873 31032
rect 279429 30680 279477 30999
rect 280813 30680 280873 30999
rect 279429 30638 280873 30680
rect 277097 26027 278517 26053
rect 277097 25773 277138 26027
rect 278478 25773 278517 26027
rect 277097 25742 278517 25773
rect 249302 19473 257654 22684
rect 250995 5327 252031 19473
rect 254084 17726 254748 17764
rect 254084 17202 254104 17726
rect 254714 17202 254748 17726
rect 254084 17150 254748 17202
rect 231680 3176 231731 4664
rect 232396 3176 232442 4664
rect 231680 582 232442 3176
rect 254084 4660 254750 17150
rect 254084 3198 254124 4660
rect 254704 3198 254750 4660
rect 254084 3110 254750 3198
rect 277273 4628 278241 25742
rect 279430 25119 280850 25144
rect 279430 24865 279469 25119
rect 280809 24865 280850 25119
rect 279430 24833 280850 24865
rect 277273 3262 277360 4628
rect 278170 3262 278241 4628
rect 277273 3177 278241 3262
rect 250995 2235 252031 2289
rect 250995 751 251034 2235
rect 251979 751 252031 2235
rect 250995 254 252031 751
rect 279693 2213 280662 24833
rect 282876 19182 283004 114932
rect 283187 91270 283510 114863
rect 283182 19182 283510 88816
rect 283688 19182 283816 114890
rect 283994 107382 284322 114862
rect 283994 32238 284322 104916
rect 284500 32238 284628 114890
rect 284806 50778 285134 114383
rect 285312 46024 285440 114890
rect 285618 46255 285946 113964
rect 286124 46024 286252 114890
rect 288812 114792 289012 115200
rect 289412 112722 289612 115349
rect 297012 114376 297212 115200
rect 297812 113954 298012 115200
rect 298212 114536 298412 115200
rect 298212 114336 298716 114536
rect 298516 112948 298716 114336
rect 286528 84302 287747 84602
rect 286528 82522 286644 84302
rect 287651 82522 287747 84302
rect 286528 4600 287747 82522
rect 286528 3247 286652 4600
rect 287645 3247 287747 4600
rect 286528 3008 287747 3247
rect 288309 80285 289528 80730
rect 288309 78505 288414 80285
rect 289421 78505 289528 80285
rect 279693 786 279768 2213
rect 280605 786 280662 2213
rect 279693 705 280662 786
rect 288309 2173 289528 78505
rect 290452 74305 291231 74519
rect 290452 69512 290546 74305
rect 291120 69512 291231 74305
rect 290452 61397 291231 69512
rect 292595 67322 293102 77663
rect 293717 74317 294224 77663
rect 293717 69482 293782 74317
rect 294150 69482 294224 74317
rect 293717 69343 294224 69482
rect 303318 74274 308118 115200
rect 311310 84307 312178 84399
rect 311310 82474 311386 84307
rect 312087 82474 312178 84307
rect 311310 77590 312178 82474
rect 311310 75481 311397 77590
rect 312080 75481 312178 77590
rect 311310 75373 312178 75481
rect 303318 69526 303458 74274
rect 308006 69526 308118 74274
rect 303318 69376 308118 69526
rect 313018 74234 317818 115200
rect 326380 113104 331160 115196
rect 336359 113104 341139 115196
rect 361812 114714 362012 115200
rect 326380 112320 341139 113104
rect 362412 112716 362612 115349
rect 385812 114228 386012 115200
rect 386412 112712 386612 115349
rect 409812 113846 410012 115200
rect 410412 112720 410612 115349
rect 433812 113410 434012 115200
rect 434412 112720 434612 115349
rect 326380 112220 331160 112320
rect 320940 93488 321264 93517
rect 319819 91499 320212 91573
rect 313018 69514 313130 74234
rect 317694 69514 317818 74234
rect 313018 69404 317818 69514
rect 315428 69400 317818 69404
rect 318960 90714 319360 90751
rect 318960 88765 319004 90714
rect 319323 88765 319360 90714
rect 292595 62487 292652 67322
rect 293020 62487 293102 67322
rect 292595 62373 293102 62487
rect 318960 67334 319360 88765
rect 319819 88736 319886 91499
rect 320160 88736 320212 91499
rect 319819 74324 320212 88736
rect 320940 91528 320963 93488
rect 321227 91528 321264 93488
rect 320940 84424 321264 91528
rect 321840 93472 322165 93500
rect 321840 91560 321890 93472
rect 322143 91560 322165 93472
rect 320940 84344 321269 84424
rect 320940 82442 320991 84344
rect 321227 82442 321269 84344
rect 320940 82378 321269 82442
rect 321840 80353 322165 91560
rect 321840 78667 321887 80353
rect 322125 78667 322165 80353
rect 326380 84230 331154 112220
rect 445288 111737 450164 115200
rect 445288 110390 445406 111737
rect 449996 110390 450164 111737
rect 445288 110133 450164 110390
rect 450478 109358 455172 115200
rect 468380 113622 473160 115224
rect 478359 113622 483139 115224
rect 503812 114296 504012 115200
rect 468380 113078 483139 113622
rect 450478 108010 450659 109358
rect 455028 108010 455172 109358
rect 450478 107772 455172 108010
rect 478359 112240 483139 113078
rect 504412 112724 504612 115349
rect 527812 114756 528012 115200
rect 528412 113118 528612 115349
rect 551812 114198 552012 115200
rect 552412 113112 552612 115349
rect 569700 114728 569900 115200
rect 570300 113124 570500 115350
rect 478359 108012 490376 112240
rect 478359 108008 483139 108012
rect 465186 106993 467270 107160
rect 354241 106521 355735 106662
rect 354241 101717 354382 106521
rect 355624 102003 355735 106521
rect 465186 105291 465393 106993
rect 467127 105291 467270 106993
rect 355624 101717 364808 102003
rect 354241 100937 364808 101717
rect 354241 100928 355735 100937
rect 352616 91801 354714 92025
rect 352616 86231 352789 91801
rect 352604 84990 352789 86231
rect 354530 84990 354714 91801
rect 352604 84786 354714 84990
rect 326380 79450 351578 84230
rect 321840 78620 322165 78667
rect 319819 69448 319884 74324
rect 320146 69448 320212 74324
rect 319819 69376 320212 69448
rect 345979 74410 346379 74420
rect 345979 74285 346385 74410
rect 345979 69476 346037 74285
rect 346312 69476 346385 74285
rect 345979 69395 346385 69476
rect 318960 62470 319016 67334
rect 319300 62470 319360 67334
rect 318960 62407 319360 62470
rect 345332 67319 345932 67433
rect 345332 62459 345399 67319
rect 345859 62459 345932 67319
rect 290452 59454 290503 61397
rect 291181 59454 291231 61397
rect 290452 27142 291231 59454
rect 345332 59110 345932 62459
rect 340532 58510 345932 59110
rect 340532 28982 341132 58510
rect 346198 58025 346385 69395
rect 346500 67296 346891 67386
rect 346500 62455 346554 67296
rect 346815 62455 346891 67296
rect 346500 62392 346891 62455
rect 342198 57838 346385 58025
rect 342198 56112 342385 57838
rect 346503 57535 346690 62392
rect 342198 55198 342211 56112
rect 342363 55198 342385 56112
rect 342198 55178 342385 55198
rect 342503 57348 346690 57535
rect 342503 56109 342690 57348
rect 342503 55217 342515 56109
rect 342664 55217 342690 56109
rect 342503 55192 342690 55217
rect 347578 53453 351578 79450
rect 352604 74295 353743 84786
rect 352604 69569 352700 74295
rect 353645 69569 353743 74295
rect 352604 69471 353743 69569
rect 352310 67250 354070 67477
rect 352310 62486 352418 67250
rect 353986 62486 354070 67250
rect 352310 59378 354070 62486
rect 352098 59225 354070 59378
rect 352098 58638 352180 59225
rect 353960 58638 354070 59225
rect 352098 58596 354070 58638
rect 352098 58578 354068 58596
rect 347578 50652 347668 53453
rect 351477 50652 351578 53453
rect 347578 50510 351578 50652
rect 339590 28602 341132 28982
rect 290452 26702 293820 27142
rect 288309 820 288423 2173
rect 289416 820 289528 2173
rect 288309 714 289528 820
rect 294461 19081 295062 19197
rect 294461 16433 294545 19081
rect 295010 16433 295062 19081
rect 294461 2206 295062 16433
rect 338710 4705 339010 18803
rect 341595 15785 341798 15803
rect 339581 15312 341096 15401
rect 339581 14892 339670 15312
rect 340952 14892 341096 15312
rect 339581 11885 341096 14892
rect 339581 11465 339692 11885
rect 340974 11465 341096 11885
rect 339581 11365 341096 11465
rect 341595 14571 341612 15785
rect 341779 14571 341798 15785
rect 338710 4669 339138 4705
rect 341595 4704 341798 14571
rect 338710 3172 338746 4669
rect 339105 3172 339138 4669
rect 338710 3133 339138 3172
rect 341465 4673 341798 4704
rect 341465 3176 341501 4673
rect 341760 3176 341798 4673
rect 341465 3142 341798 3176
rect 341595 3139 341798 3142
rect 341899 15785 342094 15806
rect 341899 14571 341910 15785
rect 342077 14571 342094 15785
rect 338712 3124 339138 3133
rect 341899 2284 342094 14571
rect 352745 14173 352885 17278
rect 342562 14033 352885 14173
rect 342562 9301 342702 14033
rect 353196 13754 353324 19139
rect 350864 13626 353324 13754
rect 353642 14328 353770 16718
rect 294461 796 294538 2206
rect 294988 796 295062 2206
rect 294461 714 295062 796
rect 341896 2237 342254 2284
rect 341896 747 341930 2237
rect 342210 747 342254 2237
rect 341896 711 342254 747
rect 346000 0 346128 7950
rect 346256 0 346384 9022
rect 346512 0 346640 7950
rect 346768 0 346896 9326
rect 347024 0 347152 7950
rect 347280 0 347408 9614
rect 347536 0 347664 7950
rect 347792 0 347920 9912
rect 348048 0 348176 7950
rect 348304 0 348432 10216
rect 348560 0 348688 7950
rect 348816 0 348944 10520
rect 349072 0 349200 7950
rect 349328 0 349456 10826
rect 349584 0 349712 7950
rect 349840 0 349968 11130
rect 350096 0 350224 7950
rect 350352 0 350480 11422
rect 350608 0 350736 7950
rect 350864 0 350992 13626
rect 353642 13325 353769 14328
rect 351376 13197 353769 13325
rect 351120 0 351248 7950
rect 351376 0 351504 13197
rect 351632 0 351760 7950
rect 351888 0 352016 10730
rect 352144 0 352272 7950
rect 352400 0 352528 11034
rect 352656 0 352784 7950
rect 352912 0 353040 11334
rect 353168 0 353296 7950
rect 353424 0 353552 11642
rect 353680 0 353808 7950
rect 353936 0 354064 11936
rect 354192 0 354320 7950
rect 354448 0 354576 12216
rect 354704 0 354832 75556
rect 354960 3114 355088 76498
rect 354960 0 355088 3068
rect 355216 0 355344 75590
rect 355472 3114 355600 76888
rect 355472 0 355600 3068
rect 355728 0 355856 75584
rect 355984 3114 356112 77304
rect 355984 0 356112 3068
rect 356240 0 356368 75578
rect 356496 3114 356624 77700
rect 356496 0 356624 3068
rect 356752 0 356880 75574
rect 357008 3114 357136 78068
rect 357008 0 357136 3068
rect 357264 0 357392 75584
rect 357520 3114 357648 78464
rect 357520 0 357648 3068
rect 357776 0 357904 75578
rect 358032 3114 358160 78860
rect 358032 0 358160 3068
rect 358288 0 358416 75564
rect 358544 3114 358672 79262
rect 358544 0 358672 3068
rect 358800 0 358928 75570
rect 359056 3114 359184 79652
rect 359056 0 359184 3068
rect 359312 0 359440 75564
rect 359568 3114 359696 80054
rect 359568 0 359696 3068
rect 359824 0 359952 75580
rect 360080 3114 360208 80450
rect 360080 0 360208 3068
rect 360336 0 360464 75578
rect 360592 3114 360720 80912
rect 360592 0 360720 3068
rect 360848 0 360976 75570
rect 361104 3114 361232 77690
rect 361104 0 361232 3068
rect 361360 0 361488 75570
rect 361616 3114 361744 77274
rect 361616 0 361744 3068
rect 361872 0 362000 75590
rect 362128 3114 362256 76878
rect 362128 0 362256 3068
rect 362384 0 362512 75590
rect 362640 3114 362768 76432
rect 362640 0 362768 3068
rect 362896 0 363024 75604
rect 363742 67288 364808 100937
rect 366265 84329 366692 84400
rect 366265 82451 366319 84329
rect 366642 82451 366692 84329
rect 366265 82391 366692 82451
rect 363742 62496 363842 67288
rect 364730 62496 364808 67288
rect 363742 62402 364808 62496
rect 365308 80389 365509 80395
rect 365308 80321 365736 80389
rect 365308 78476 365384 80321
rect 365659 78476 365736 80321
rect 365308 78390 365736 78476
rect 365870 80311 366207 80395
rect 365870 78432 365904 80311
rect 366152 78432 366207 80311
rect 365308 61754 365509 78390
rect 365870 78188 366207 78432
rect 364735 61553 365509 61754
rect 364735 50211 364936 61553
rect 364735 49357 364765 50211
rect 364915 49357 364936 50211
rect 364735 49322 364936 49357
rect 366450 49435 366692 82391
rect 366966 84346 367303 84393
rect 366966 82450 367001 84346
rect 367267 82450 367303 84346
rect 366966 78187 367303 82450
rect 371592 84346 371929 84393
rect 371592 82450 371627 84346
rect 371893 82450 371929 84346
rect 370496 80311 370832 80395
rect 370496 78432 370530 80311
rect 370778 78432 370832 80311
rect 370496 78188 370832 78432
rect 371592 78187 371929 82450
rect 374682 84318 375243 84392
rect 374682 82435 374726 84318
rect 375181 82435 375243 84318
rect 374682 79563 375243 82435
rect 376218 84346 376555 84393
rect 376218 82450 376253 84346
rect 376519 82450 376555 84346
rect 374682 79434 374700 79563
rect 375223 79434 375243 79563
rect 374682 79411 375243 79434
rect 375477 80350 376122 80389
rect 375477 80126 375516 80350
rect 376086 80126 376122 80350
rect 375477 79999 375497 80126
rect 376097 79999 376122 80126
rect 375477 78889 375516 79999
rect 375440 78432 375516 78889
rect 376086 78432 376122 79999
rect 375440 78392 376122 78432
rect 368214 74363 368551 77843
rect 368214 69414 368232 74363
rect 368531 69414 368551 74363
rect 368214 69387 368551 69414
rect 369838 67349 370175 77845
rect 372840 74363 373177 77840
rect 374464 76749 374801 77836
rect 375440 77821 375755 78392
rect 376218 78187 376555 82450
rect 380844 84346 381181 84393
rect 380844 82450 380879 84346
rect 381145 82450 381181 84346
rect 373462 76744 374801 76749
rect 372840 69414 372858 74363
rect 373157 69414 373177 74363
rect 372840 69387 373177 69414
rect 373461 76412 374801 76744
rect 373461 67417 373888 76412
rect 369838 62448 369876 67349
rect 370126 62448 370175 67349
rect 369838 62407 370175 62448
rect 372250 67295 373888 67417
rect 372250 62506 372355 67295
rect 373406 65842 373888 67295
rect 374299 74290 375345 74424
rect 374299 69477 374411 74290
rect 375214 69477 375345 74290
rect 373406 62506 373523 65842
rect 372250 59420 373523 62506
rect 372250 58463 372341 59420
rect 373424 58463 373523 59420
rect 372250 58359 373523 58463
rect 374299 52920 375345 69477
rect 374299 52579 374345 52920
rect 375302 52579 375345 52920
rect 374299 52526 375345 52579
rect 376007 74328 376909 74425
rect 376007 69459 376090 74328
rect 376822 69459 376909 74328
rect 366450 49395 369247 49435
rect 366450 49227 368319 49395
rect 369200 49227 369247 49395
rect 366450 49193 369247 49227
rect 376007 48638 376909 69459
rect 377466 74363 377803 80946
rect 377466 69414 377484 74363
rect 377783 69414 377803 74363
rect 377466 69387 377803 69414
rect 364508 47736 376909 48638
rect 378099 67323 379001 67430
rect 378099 62448 378163 67323
rect 378932 62448 379001 67323
rect 363174 21284 363548 21318
rect 363174 20548 363198 21284
rect 363516 20548 363548 21284
rect 363174 20524 363548 20548
rect 363174 6930 363278 20524
rect 364508 16947 365410 47736
rect 378099 47278 379001 62448
rect 379090 67349 379427 82418
rect 379948 80311 380284 80395
rect 379948 78432 379982 80311
rect 380230 78432 380284 80311
rect 379948 78188 380284 78432
rect 380844 78187 381181 82450
rect 385422 84350 386120 84411
rect 385422 82438 385474 84350
rect 386053 82438 386120 84350
rect 384374 80394 384710 80395
rect 384357 80337 385102 80394
rect 384357 78432 384408 80337
rect 385036 78432 385102 80337
rect 382092 74363 382429 77840
rect 382092 69414 382110 74363
rect 382409 69414 382429 74363
rect 382092 69387 382429 69414
rect 379090 62448 379128 67349
rect 379378 62448 379427 67349
rect 379090 62407 379427 62448
rect 383716 67349 384053 77843
rect 383716 62448 383754 67349
rect 384004 62448 384053 67349
rect 383716 62407 384053 62448
rect 382912 53463 383955 53537
rect 382912 50614 382998 53463
rect 383893 50614 383955 53463
rect 382912 50530 383955 50614
rect 364508 15024 364589 16947
rect 365295 15024 365410 16947
rect 364508 14949 365410 15024
rect 365743 46376 379001 47278
rect 365743 16970 366645 46376
rect 368182 45515 369817 45667
rect 368182 45451 368294 45515
rect 368180 44750 368294 45451
rect 369665 44750 369817 45515
rect 368180 44591 369817 44750
rect 368180 43841 368577 44591
rect 383168 39215 383713 50530
rect 384357 41662 385102 78432
rect 385422 43750 386120 82438
rect 388876 84328 389391 89266
rect 388876 82465 388948 84328
rect 389318 82843 389391 84328
rect 389318 82465 389695 82843
rect 388876 82404 389695 82465
rect 388876 82403 389391 82404
rect 389000 80311 389336 80395
rect 389000 78432 389034 80311
rect 389282 78432 389336 80311
rect 389000 78188 389336 78432
rect 389469 78190 389695 82404
rect 389830 80315 390448 90955
rect 389830 78524 389905 80315
rect 390347 78524 390448 80315
rect 389830 78416 390448 78524
rect 389469 77964 390101 78190
rect 386718 74363 387055 77840
rect 386718 69414 386736 74363
rect 387035 69414 387055 74363
rect 386718 69387 387055 69414
rect 388342 67349 388679 77843
rect 390853 76243 390993 92951
rect 388342 62448 388380 67349
rect 388630 62448 388679 67349
rect 388342 62407 388679 62448
rect 388839 76103 390993 76243
rect 385241 43716 386120 43750
rect 385241 43242 385274 43716
rect 386087 43242 386120 43716
rect 385241 43227 386120 43242
rect 385241 43211 386119 43227
rect 384012 41614 385956 41662
rect 384012 41169 384078 41614
rect 385891 41169 385956 41614
rect 384012 41112 385956 41169
rect 372113 38670 383713 39215
rect 384352 39680 385786 39728
rect 384352 39126 384400 39680
rect 385734 39126 385786 39680
rect 384352 39078 385786 39126
rect 386280 18518 386406 61225
rect 387016 19536 387153 60358
rect 387733 21120 387877 61577
rect 388394 20215 388531 61871
rect 388839 19812 388979 76103
rect 391353 73672 391493 94425
rect 391654 74343 391988 77839
rect 391654 69422 391692 74343
rect 391938 69422 391988 74343
rect 392053 73152 392193 95726
rect 399348 84346 399685 84393
rect 403974 84392 404311 84393
rect 395335 84285 395702 84316
rect 393939 83338 394612 83416
rect 392403 75381 392650 77847
rect 392856 76317 393476 81258
rect 393939 80729 394019 83338
rect 394553 80729 394612 83338
rect 393939 79820 394612 80729
rect 394806 82606 395189 82668
rect 394806 80687 394851 82606
rect 395147 80687 395189 82606
rect 394806 80393 395189 80687
rect 395335 82442 395377 84285
rect 395670 82442 395702 84285
rect 395335 81521 395702 82442
rect 399348 82450 399383 84346
rect 399649 82450 399685 84346
rect 395335 81462 395710 81521
rect 395335 80671 395370 81462
rect 395671 80936 395710 81462
rect 395671 80671 395711 80936
rect 395335 80626 395711 80671
rect 394806 80338 395289 80393
rect 394806 80044 394948 80338
rect 393939 79108 394692 79820
rect 393559 78889 393907 78943
rect 393559 78434 393607 78889
rect 393862 78434 393907 78889
rect 393559 77831 393907 78434
rect 394019 77323 394692 79108
rect 394906 78459 394948 80044
rect 395252 78459 395289 80338
rect 394906 78391 395289 78459
rect 395437 78200 395711 80626
rect 395118 77926 395711 78200
rect 396646 80346 397300 80416
rect 396646 78431 396692 80346
rect 397253 78431 397300 80346
rect 394019 76650 395320 77323
rect 392856 75697 394280 76317
rect 392403 75134 393458 75381
rect 391654 69372 391988 69422
rect 393211 67400 393458 75134
rect 393660 74321 394280 75697
rect 393660 69498 393729 74321
rect 394202 69498 394280 74321
rect 393660 69405 394280 69498
rect 393210 67327 393598 67400
rect 393210 62461 393277 67327
rect 393531 62461 393598 67327
rect 393210 62388 393598 62461
rect 394647 67323 395320 76650
rect 395970 74363 396307 77840
rect 395970 69414 395988 74363
rect 396287 69414 396307 74363
rect 395970 69387 396307 69414
rect 394647 62485 394738 67323
rect 395227 62485 395320 67323
rect 394647 62404 395320 62485
rect 396646 60288 397300 78431
rect 398252 80311 398588 80395
rect 398252 78432 398286 80311
rect 398534 78432 398588 80311
rect 398252 78188 398588 78432
rect 399348 78187 399685 82450
rect 403760 84347 404313 84392
rect 403760 82436 403823 84347
rect 404281 82436 404313 84347
rect 402878 80341 403417 80403
rect 402878 78432 402912 80341
rect 403367 78432 403417 80341
rect 397594 67349 397931 77843
rect 400596 74363 400933 77840
rect 400596 69414 400614 74363
rect 400913 69414 400933 74363
rect 400596 69387 400933 69414
rect 397594 62448 397632 67349
rect 397882 62448 397931 67349
rect 397594 62407 397931 62448
rect 402220 67349 402557 77843
rect 402220 62448 402258 67349
rect 402508 62448 402557 67349
rect 402220 62407 402557 62448
rect 402878 60612 403417 78432
rect 393128 59634 397300 60288
rect 399435 60073 403417 60612
rect 403760 60624 404313 82436
rect 408600 84346 408937 84393
rect 408600 82450 408635 84346
rect 408901 82450 408937 84346
rect 407504 80311 407840 80395
rect 407504 78432 407538 80311
rect 407786 78432 407840 80311
rect 407504 78188 407840 78432
rect 408600 78187 408937 82450
rect 413226 84346 413563 84393
rect 413226 82450 413261 84346
rect 413527 82450 413563 84346
rect 412130 80311 412466 80395
rect 412130 78432 412164 80311
rect 412412 78432 412466 80311
rect 412130 78188 412466 78432
rect 413226 78187 413563 82450
rect 417852 84346 418189 84393
rect 417852 82450 417887 84346
rect 418153 82450 418189 84346
rect 416756 80311 417092 80395
rect 416756 78432 416790 80311
rect 417038 78432 417092 80311
rect 416756 78188 417092 78432
rect 417852 78187 418189 82450
rect 422478 84346 422815 84393
rect 422478 82450 422513 84346
rect 422779 82450 422815 84346
rect 421382 80311 421718 80395
rect 421382 78432 421416 80311
rect 421664 78432 421718 80311
rect 421382 78188 421718 78432
rect 422478 78187 422815 82450
rect 424314 84339 424642 84381
rect 424314 82430 424351 84339
rect 424599 82430 424642 84339
rect 431730 84346 432067 84393
rect 405222 74363 405559 77840
rect 405222 69414 405240 74363
rect 405539 69414 405559 74363
rect 405222 69387 405559 69414
rect 406846 67349 407183 77843
rect 409848 74363 410185 77840
rect 409848 69414 409866 74363
rect 410165 69414 410185 74363
rect 409848 69387 410185 69414
rect 406846 62448 406884 67349
rect 407134 62448 407183 67349
rect 406846 62407 407183 62448
rect 411472 67349 411809 77843
rect 414474 74363 414811 77840
rect 414474 69414 414492 74363
rect 414791 69414 414811 74363
rect 414474 69387 414811 69414
rect 411472 62448 411510 67349
rect 411760 62448 411809 67349
rect 411472 62407 411809 62448
rect 416098 67349 416435 77843
rect 419100 74363 419437 77840
rect 419100 69414 419118 74363
rect 419417 69414 419437 74363
rect 419100 69387 419437 69414
rect 416098 62448 416136 67349
rect 416386 62448 416435 67349
rect 416098 62407 416435 62448
rect 420724 67349 421061 77843
rect 422518 74339 423268 74433
rect 422518 69456 422587 74339
rect 423195 69456 423268 74339
rect 420724 62448 420762 67349
rect 421012 62448 421061 67349
rect 420724 62407 421061 62448
rect 421472 67324 422241 67410
rect 421472 62471 421550 67324
rect 422153 62471 422241 67324
rect 414838 61829 415704 61941
rect 414838 60678 414932 61829
rect 415612 60678 415704 61829
rect 389684 53468 391062 53564
rect 389684 50582 389744 53468
rect 390995 50582 391062 53468
rect 389684 32738 391062 50582
rect 389684 32467 389701 32738
rect 391045 32467 391062 32738
rect 389684 32431 391062 32467
rect 391399 48413 392808 48502
rect 391399 45614 391494 48413
rect 392733 45614 392808 48413
rect 391399 29129 392808 45614
rect 393134 31332 393549 59634
rect 399435 53451 399974 60073
rect 403760 60071 405080 60624
rect 414838 60575 415704 60678
rect 421472 60080 422241 62471
rect 404527 53483 405080 60071
rect 405417 59916 406547 59944
rect 405417 59616 405465 59916
rect 406501 59616 406547 59916
rect 405417 59583 406547 59616
rect 399435 52912 403417 53451
rect 402878 45342 403417 52912
rect 402878 44613 402922 45342
rect 403374 44613 403417 45342
rect 403760 52930 405080 53483
rect 403760 45940 404313 52930
rect 403760 44919 403806 45940
rect 404042 44919 404313 45940
rect 405446 48473 406518 59583
rect 414900 59311 422241 60080
rect 422518 60764 423268 69456
rect 423726 74363 424063 77840
rect 423726 69414 423744 74363
rect 424043 69414 424063 74363
rect 423726 69387 424063 69414
rect 424314 61455 424642 82430
rect 427349 84189 427741 84235
rect 427349 82476 427404 84189
rect 427681 82476 427741 84189
rect 428452 83660 429116 83735
rect 427349 81455 427741 82476
rect 427887 82532 428289 82602
rect 427342 81409 427744 81455
rect 427342 80985 427385 81409
rect 427104 80611 427385 80985
rect 427699 80611 427744 81409
rect 427104 80571 427744 80611
rect 427887 80638 427915 82532
rect 428234 80638 428289 82532
rect 424787 80347 425115 80418
rect 424787 78438 424822 80347
rect 425070 78438 425115 80347
rect 424787 62029 425115 78438
rect 426008 80311 426344 80395
rect 426008 78432 426042 80311
rect 426290 78432 426344 80311
rect 426008 78188 426344 78432
rect 427104 78195 427441 80571
rect 427887 80342 428289 80638
rect 427887 78463 427942 80342
rect 428243 78463 428289 80342
rect 427887 78392 428289 78463
rect 428452 80656 428533 83660
rect 429062 80656 429116 83660
rect 431730 82450 431765 84346
rect 432031 82450 432067 84346
rect 425350 67349 425687 77843
rect 427952 74338 428289 77849
rect 427952 69455 427997 74338
rect 428235 69455 428289 74338
rect 427952 69404 428289 69455
rect 425350 62448 425388 67349
rect 425638 62448 425687 67349
rect 425350 62407 425687 62448
rect 428452 67316 429116 80656
rect 429480 74290 430100 81198
rect 430934 80311 431270 80395
rect 430934 78432 430968 80311
rect 431216 78432 431270 80311
rect 430934 78188 431270 78432
rect 431730 78187 432067 82450
rect 429480 69452 429574 74290
rect 430005 69452 430100 74290
rect 429480 69373 430100 69452
rect 428452 62479 428531 67316
rect 429041 62479 429116 67316
rect 428452 62381 429116 62479
rect 430276 67349 430613 77841
rect 432359 74162 432499 95756
rect 432859 74683 432999 94455
rect 433159 75361 433496 77847
rect 433659 76235 433799 92981
rect 434234 80333 434813 90809
rect 435229 84337 435807 89282
rect 435229 82453 435287 84337
rect 435737 82453 435807 84337
rect 435229 82378 435807 82453
rect 436356 84346 436693 84393
rect 436356 82450 436391 84346
rect 436657 82450 436693 84346
rect 434234 78449 434297 80333
rect 434747 78449 434813 80333
rect 434234 78388 434813 78449
rect 435260 80311 435596 80395
rect 435260 78432 435294 80311
rect 435542 78432 435596 80311
rect 435260 78188 435596 78432
rect 436356 78187 436693 82450
rect 440982 84346 441319 84393
rect 440982 82450 441017 84346
rect 441283 82450 441319 84346
rect 440056 80311 440392 80395
rect 440056 78432 440090 80311
rect 440338 78432 440392 80311
rect 440056 78188 440392 78432
rect 440982 78187 441319 82450
rect 445608 84346 445945 84393
rect 445608 82450 445643 84346
rect 445909 82450 445945 84346
rect 444682 80311 445018 80395
rect 444682 78432 444716 80311
rect 444964 78432 445018 80311
rect 444682 78188 445018 78432
rect 445608 78187 445945 82450
rect 450234 84346 450571 84393
rect 450234 82450 450269 84346
rect 450535 82450 450571 84346
rect 449138 80311 449474 80395
rect 449138 78432 449172 80311
rect 449420 78432 449474 80311
rect 449138 78188 449474 78432
rect 450234 78187 450571 82450
rect 451647 84338 452298 84397
rect 451647 82445 451692 84338
rect 452265 82445 452298 84338
rect 454860 84346 455197 84393
rect 450732 80358 451400 80400
rect 450732 80303 450780 80358
rect 451361 80303 451400 80358
rect 450732 80161 450757 80303
rect 451373 80161 451400 80303
rect 450732 78430 450780 80161
rect 451361 78430 451400 80161
rect 451647 79631 452298 82445
rect 451647 79499 451681 79631
rect 452277 79499 452298 79631
rect 451647 79469 452298 79499
rect 450732 78382 451400 78430
rect 434602 76890 434939 77836
rect 434602 76553 435400 76890
rect 433659 76095 434833 76235
rect 433159 75024 434328 75361
rect 433991 74329 434328 75024
rect 433991 70845 434031 74329
rect 434276 70845 434328 74329
rect 433991 70786 434328 70845
rect 434693 70583 434833 76095
rect 430276 62443 430327 67349
rect 430568 62443 430613 67349
rect 430276 62371 430613 62443
rect 430906 70443 434833 70583
rect 424787 61701 430665 62029
rect 424314 61127 430192 61455
rect 422518 60014 429638 60764
rect 414900 52381 415669 59311
rect 414900 51919 422027 52381
rect 414900 51773 421070 51919
rect 421767 51773 422027 51919
rect 414900 51612 422027 51773
rect 428888 50307 429638 60014
rect 421022 49557 429638 50307
rect 421022 48515 421772 49557
rect 405446 45583 405504 48473
rect 406457 45583 406518 48473
rect 421004 48487 421774 48515
rect 421004 48341 421046 48487
rect 421743 48341 421774 48487
rect 421004 48310 421774 48341
rect 429864 47261 430192 61127
rect 420743 47148 430192 47261
rect 420743 47023 420803 47148
rect 421743 47023 430192 47148
rect 420743 46933 430192 47023
rect 430337 46281 430665 61701
rect 420728 46173 430665 46281
rect 420728 46034 420789 46173
rect 421670 46034 430665 46173
rect 420728 45953 430665 46034
rect 405446 45522 406518 45583
rect 403760 44879 404313 44919
rect 402878 44550 403417 44613
rect 391399 29084 393015 29129
rect 391399 28593 391451 29084
rect 392975 28593 393015 29084
rect 391399 28566 393015 28593
rect 391405 28550 393015 28566
rect 430906 20798 431046 70443
rect 431401 67324 432219 67472
rect 431401 62472 431483 67324
rect 432140 62472 432219 67324
rect 431401 22898 432219 62472
rect 435063 67346 435400 76553
rect 437604 74363 437941 77840
rect 437604 69414 437622 74363
rect 437921 69414 437941 74363
rect 437604 69387 437941 69414
rect 435063 62462 435109 67346
rect 435349 62462 435400 67346
rect 435063 62398 435400 62462
rect 439228 67349 439565 77843
rect 442230 74363 442567 77840
rect 442230 69414 442248 74363
rect 442547 69414 442567 74363
rect 442230 69387 442567 69414
rect 439228 62448 439266 67349
rect 439516 62448 439565 67349
rect 439228 62407 439565 62448
rect 443854 67349 444191 77843
rect 446856 74363 447193 77840
rect 446856 69414 446874 74363
rect 447173 69414 447193 74363
rect 446856 69387 447193 69414
rect 443854 62448 443892 67349
rect 444142 62448 444191 67349
rect 443854 62407 444191 62448
rect 448480 67349 448817 77843
rect 451482 74363 451819 77840
rect 451482 69414 451500 74363
rect 451799 69414 451819 74363
rect 451482 69387 451819 69414
rect 448480 62448 448518 67349
rect 448768 62448 448817 67349
rect 448480 62407 448817 62448
rect 453006 67349 453343 82514
rect 454860 82450 454895 84346
rect 455161 82450 455197 84346
rect 453934 80311 454270 80395
rect 453934 78432 453968 80311
rect 454216 78432 454270 80311
rect 453934 78188 454270 78432
rect 454860 78187 455197 82450
rect 459486 84346 459823 84393
rect 459486 82450 459521 84346
rect 459787 82450 459823 84346
rect 456108 74363 456445 81110
rect 458590 80311 458926 80395
rect 458590 78432 458624 80311
rect 458872 78432 458926 80311
rect 458590 78188 458926 78432
rect 459486 78187 459823 82450
rect 464112 84346 464449 84393
rect 464112 82450 464147 84346
rect 464413 82450 464449 84346
rect 463116 80311 463452 80395
rect 463116 78432 463150 80311
rect 463398 78432 463452 80311
rect 463116 78188 463452 78432
rect 464112 78187 464449 82450
rect 456108 69414 456126 74363
rect 456425 69414 456445 74363
rect 456108 69387 456445 69414
rect 453006 62448 453044 67349
rect 453294 62448 453343 67349
rect 453006 62407 453343 62448
rect 457732 67349 458069 77843
rect 460734 74363 461071 77840
rect 460734 69414 460752 74363
rect 461051 69414 461071 74363
rect 460734 69387 461071 69414
rect 457732 62448 457770 67349
rect 458020 62448 458069 67349
rect 457732 62407 458069 62448
rect 462158 67349 462495 77843
rect 464660 74342 464997 77842
rect 464660 69463 464711 74342
rect 464949 69463 464997 74342
rect 464660 69399 464997 69463
rect 462158 62448 462196 67349
rect 462446 62448 462495 67349
rect 462158 62407 462495 62448
rect 465186 67277 467270 105291
rect 486148 89522 490376 108012
rect 508078 110004 508814 110093
rect 508078 109535 508087 110004
rect 508795 109535 508814 110004
rect 473606 86252 475524 86410
rect 473606 84830 473636 86252
rect 475432 85748 475524 86252
rect 486148 86228 486280 89522
rect 490240 86228 490376 89522
rect 486148 86098 490376 86228
rect 475432 84830 475957 85748
rect 473606 84754 475957 84830
rect 468738 84346 469075 84393
rect 468738 82450 468773 84346
rect 469039 82450 469075 84346
rect 467842 80311 468178 80395
rect 467842 78432 467876 80311
rect 468124 78432 468178 80311
rect 467842 78188 468178 78432
rect 468738 78187 469075 82450
rect 473364 84346 473701 84393
rect 473364 82450 473399 84346
rect 473665 82450 473701 84346
rect 472468 80311 472804 80395
rect 472468 78432 472502 80311
rect 472750 78432 472804 80311
rect 472468 78188 472804 78432
rect 473364 78187 473701 82450
rect 469986 74363 470323 77840
rect 469986 69414 470004 74363
rect 470303 69414 470323 74363
rect 469986 69387 470323 69414
rect 465186 62510 465312 67277
rect 467131 62510 467270 67277
rect 465186 62268 467270 62510
rect 471210 67349 471547 77843
rect 473911 74237 475957 84754
rect 484883 85112 489190 85252
rect 477949 84346 478802 84425
rect 477949 82450 478025 84346
rect 478291 84345 478802 84346
rect 478720 82450 478802 84345
rect 477094 80391 477430 80395
rect 476762 80342 477619 80391
rect 476762 78423 476801 80342
rect 477563 78423 477619 80342
rect 473911 69572 474098 74237
rect 475813 69572 475957 74237
rect 473911 69406 475957 69572
rect 471210 62448 471248 67349
rect 471498 62448 471547 67349
rect 471210 62407 471547 62448
rect 476136 67349 476473 77843
rect 476136 62448 476174 67349
rect 476424 62448 476473 67349
rect 476136 62407 476473 62448
rect 476762 59794 477619 78423
rect 477949 59826 478802 82450
rect 482616 84346 482953 84393
rect 482616 82450 482651 84346
rect 482917 82450 482953 84346
rect 481720 80311 482056 80395
rect 481720 78432 481754 80311
rect 482002 78432 482056 80311
rect 481720 78188 482056 78432
rect 482616 78187 482953 82450
rect 479238 74363 479575 77840
rect 479238 69414 479256 74363
rect 479555 69414 479575 74363
rect 479238 69387 479575 69414
rect 480862 67349 481199 77843
rect 483864 74409 484201 77852
rect 484883 75522 485023 85112
rect 491214 85012 491374 99052
rect 489734 84852 491374 85012
rect 487242 84346 487579 84393
rect 487242 82450 487277 84346
rect 487543 82450 487579 84346
rect 486346 80311 486682 80395
rect 486346 78432 486380 80311
rect 486628 78432 486682 80311
rect 486346 78188 486682 78432
rect 487242 78187 487579 82450
rect 485388 76580 485725 77841
rect 485388 76243 486586 76580
rect 484883 75382 486050 75522
rect 483864 74249 485626 74409
rect 483864 74004 484043 74249
rect 480862 62448 480900 67349
rect 481150 62448 481199 67349
rect 483909 69527 484043 74004
rect 485525 69527 485626 74249
rect 483909 64842 485626 69527
rect 480862 62407 481199 62448
rect 482509 63142 485626 64842
rect 473864 58834 477619 59794
rect 474592 55184 475929 55264
rect 477901 45966 478861 59826
rect 432479 31895 433187 45918
rect 474624 45006 478861 45966
rect 482509 43514 484226 63142
rect 485910 62547 486050 75382
rect 484636 62407 486050 62547
rect 486249 67394 486586 76243
rect 488490 74433 488827 77852
rect 489734 77454 489894 84852
rect 492652 84712 492812 106882
rect 498225 93854 498552 93932
rect 498225 91530 498275 93854
rect 498510 91530 498552 93854
rect 491436 84552 492814 84712
rect 490972 80311 491308 80395
rect 490972 78432 491006 80311
rect 491254 78432 491308 80311
rect 490972 78188 491308 78432
rect 490114 75617 490451 77844
rect 491436 77058 491596 84552
rect 491868 84346 492205 84393
rect 491868 82450 491903 84346
rect 492169 82450 492205 84346
rect 491868 78187 492205 82450
rect 496494 84346 496831 84393
rect 496494 82450 496529 84346
rect 496795 82450 496831 84346
rect 495598 80311 495934 80395
rect 495598 78432 495632 80311
rect 495880 78432 495934 80311
rect 495598 78188 495934 78432
rect 496494 78187 496831 82450
rect 498225 80325 498552 91530
rect 499144 93829 499471 93932
rect 499144 91505 499190 93829
rect 499425 91505 499471 93829
rect 499144 84409 499471 91505
rect 504041 93849 504432 93904
rect 504041 91513 504104 93849
rect 504385 91513 504432 93849
rect 499144 84323 499511 84409
rect 499144 82442 499199 84323
rect 499453 82442 499511 84323
rect 501120 84346 501457 84393
rect 499144 82386 499511 82442
rect 499924 84146 500260 84180
rect 499924 82893 499949 84146
rect 500235 82893 500260 84146
rect 498225 78443 498269 80325
rect 498514 78443 498552 80325
rect 498225 78361 498552 78443
rect 499924 80311 500260 82893
rect 499924 78432 499958 80311
rect 500206 78432 500260 80311
rect 499924 78188 500260 78432
rect 501120 83150 501155 84346
rect 501120 81984 501152 83150
rect 501421 82450 501457 84346
rect 504041 82672 504432 91513
rect 501407 81984 501457 82450
rect 501120 78187 501457 81984
rect 502348 82281 504432 82672
rect 505066 93832 505457 93904
rect 505066 91496 505121 93832
rect 505402 91496 505457 93832
rect 490114 75280 491137 75617
rect 488490 74302 490404 74433
rect 488490 74004 488817 74302
rect 488719 69518 488817 74004
rect 490270 69518 490404 74302
rect 486249 67310 486626 67394
rect 486249 62481 486318 67310
rect 486562 62481 486626 67310
rect 482509 43140 484224 43514
rect 432479 31571 432505 31895
rect 433161 31571 433187 31895
rect 432479 31545 433187 31571
rect 431401 22716 434989 22898
rect 431401 21830 432014 22716
rect 434717 21830 434989 22716
rect 431401 21558 434989 21830
rect 435460 19028 435614 42893
rect 451984 42872 484224 43140
rect 451984 41819 452319 42872
rect 459350 41819 484224 42872
rect 451984 41551 484224 41819
rect 484636 40403 484776 62407
rect 486249 62401 486626 62481
rect 486883 67294 488568 67398
rect 486883 62510 487006 67294
rect 488459 62510 488568 67294
rect 486883 59935 488568 62510
rect 488719 59969 490404 69518
rect 490800 67346 491137 75280
rect 493116 74363 493453 77840
rect 493116 69414 493134 74363
rect 493433 69414 493453 74363
rect 493116 69387 493453 69414
rect 490800 62471 490841 67346
rect 491077 62471 491137 67346
rect 490800 62400 491137 62471
rect 494540 67349 494877 77843
rect 497742 74404 498079 77849
rect 499366 75610 499703 77841
rect 502348 77261 502739 82281
rect 505066 81852 505457 91496
rect 504008 81461 505457 81852
rect 504008 77843 504399 81461
rect 503992 77359 504399 77843
rect 499366 75273 500701 75610
rect 494540 62448 494578 67349
rect 494828 62448 494877 67349
rect 494540 62407 494877 62448
rect 496423 74294 498108 74404
rect 496423 69510 496534 74294
rect 497987 69510 498108 74294
rect 496423 59967 498108 69510
rect 498259 67291 499944 67390
rect 498259 62507 498357 67291
rect 499810 62507 499944 67291
rect 498259 59980 499944 62507
rect 500364 67353 500701 75273
rect 502368 74363 502705 77261
rect 502368 69414 502386 74363
rect 502685 69414 502705 74363
rect 502368 69387 502705 69414
rect 503992 67690 504329 77359
rect 505854 76674 506014 106560
rect 506672 76252 506832 98692
rect 508078 82112 508814 109535
rect 508078 81348 508114 82112
rect 508775 81348 508814 82112
rect 508078 74444 508814 81348
rect 509036 108138 509652 108159
rect 509036 107636 509061 108138
rect 509627 107636 509652 108138
rect 509036 83514 509652 107636
rect 573656 95095 573956 95105
rect 554170 89337 555098 89376
rect 509036 82928 509068 83514
rect 509620 82928 509652 83514
rect 500364 62445 500401 67353
rect 500662 62445 500701 67353
rect 500364 62393 500701 62445
rect 503742 67361 504329 67690
rect 507199 74313 508884 74444
rect 507199 69529 507329 74313
rect 508782 69529 508884 74313
rect 503742 67349 504079 67361
rect 503742 62448 503780 67349
rect 504030 62448 504079 67349
rect 503742 62407 504079 62448
rect 505363 67262 507048 67398
rect 505363 62478 505496 67262
rect 506949 62478 507048 67262
rect 505363 59935 507048 62478
rect 507199 59980 508884 69529
rect 509036 67391 509652 82928
rect 511039 89021 515267 89201
rect 511039 85727 511154 89021
rect 515114 85727 515267 89021
rect 554170 89107 554213 89337
rect 555054 89107 555098 89337
rect 511039 80662 515267 85727
rect 552681 88427 553924 88460
rect 552681 88193 552725 88427
rect 553869 88193 553924 88427
rect 535535 84427 535855 84430
rect 535385 84314 535855 84427
rect 532826 83634 533280 83671
rect 532826 82455 532883 83634
rect 533201 82455 533280 83634
rect 511039 76434 525562 80662
rect 514908 74294 516593 74404
rect 514908 69510 515008 74294
rect 516461 69510 516593 74294
rect 509021 67281 510709 67391
rect 509021 66694 509143 67281
rect 509024 62497 509143 66694
rect 510596 62497 510709 67281
rect 509024 62384 510709 62497
rect 509036 62193 509652 62384
rect 514908 59999 516593 69510
rect 516741 67281 518429 67391
rect 516741 66694 516863 67281
rect 516744 62497 516863 66694
rect 518316 62497 518429 67281
rect 516744 59990 518429 62497
rect 521334 48410 525562 76434
rect 526663 63960 526915 79767
rect 530546 74316 530945 74433
rect 530546 69458 530609 74316
rect 530860 69458 530945 74316
rect 529537 67324 529936 67406
rect 529537 62466 529618 67324
rect 529869 62466 529936 67324
rect 521334 45689 521477 48410
rect 525395 45689 525562 48410
rect 521334 45518 525562 45689
rect 483337 40263 484776 40403
rect 479068 38784 480580 38984
rect 479068 34694 479268 38784
rect 480424 34694 480580 38784
rect 472975 22662 478554 22814
rect 472975 21637 473177 22662
rect 478353 21637 478554 22662
rect 472975 21503 478554 21637
rect 475586 19501 478387 21503
rect 452216 19330 463985 19470
rect 441122 18850 453924 18990
rect 441122 17304 441262 18850
rect 463831 18029 463971 19330
rect 479068 20475 480580 34694
rect 479068 18553 479182 20475
rect 480378 18553 480580 20475
rect 479068 18337 480580 18553
rect 483337 18029 483477 40263
rect 463831 17889 483477 18029
rect 461239 17462 484333 17601
rect 415459 17164 441262 17304
rect 365743 15047 365875 16970
rect 366581 15047 366645 16970
rect 416265 16561 429536 16728
rect 429369 16286 429536 16561
rect 467449 16552 483869 16729
rect 429369 16119 438791 16286
rect 464295 15163 483528 15317
rect 365743 14966 366645 15047
rect 364534 2226 365054 9425
rect 485124 9393 486684 12274
rect 487522 10794 488298 10844
rect 487522 10414 487572 10794
rect 488240 10414 488298 10794
rect 487522 10356 488298 10414
rect 482997 8193 486684 9393
rect 475454 7697 476850 7849
rect 457691 7228 458056 7291
rect 457691 6898 457704 7228
rect 458043 6898 458056 7228
rect 457691 6530 458056 6898
rect 468366 7245 468731 7264
rect 468366 6914 468381 7245
rect 468715 6914 468731 7245
rect 468366 6530 468731 6914
rect 457691 6165 468731 6530
rect 475454 6385 475597 7697
rect 476706 6385 476850 7697
rect 364534 770 364588 2226
rect 365003 770 365054 2226
rect 364534 704 365054 770
rect 475454 2136 476850 6385
rect 475454 824 475597 2136
rect 476706 824 476850 2136
rect 475454 723 476850 824
rect 485124 2202 486684 8193
rect 490606 4624 492006 12295
rect 490606 3276 490718 4624
rect 491898 3276 492006 4624
rect 490606 3020 492006 3276
rect 494836 4638 496088 10972
rect 494836 3202 494902 4638
rect 496002 3202 496088 4638
rect 494836 3100 496088 3202
rect 485124 843 485221 2202
rect 486580 843 486684 2202
rect 485124 616 486684 843
rect 500236 2210 501433 10994
rect 500236 774 500288 2210
rect 501388 774 501433 2210
rect 500236 702 501433 774
rect 503844 2172 505084 11103
rect 509240 4588 510458 11136
rect 509240 3217 509316 4588
rect 510361 3217 510458 4588
rect 509240 3119 510458 3217
rect 513355 4634 514555 10322
rect 513355 3198 513408 4634
rect 514508 3198 514555 4634
rect 513355 3100 514555 3198
rect 503844 801 503942 2172
rect 504987 801 505084 2172
rect 503844 693 505084 801
rect 518727 2210 519927 10234
rect 526602 7794 526812 61949
rect 527130 34314 527350 60712
rect 527668 47690 527888 60540
rect 529537 58947 529936 62466
rect 529537 57678 529578 58947
rect 529863 57678 529936 58947
rect 529537 57604 529936 57678
rect 530546 58995 530945 69458
rect 530546 57726 530611 58995
rect 530896 57726 530945 58995
rect 530546 57637 530945 57726
rect 528152 9050 528431 33492
rect 530704 15879 530969 47415
rect 532826 41065 533280 82455
rect 535385 82458 535463 84314
rect 535798 82458 535855 84314
rect 535385 82391 535855 82458
rect 532826 40806 532870 41065
rect 533236 40806 533280 41065
rect 531331 16331 531596 34140
rect 532826 27508 533280 40806
rect 532826 27232 532860 27508
rect 533256 27232 533280 27508
rect 532826 21069 533280 27232
rect 533674 80331 534128 80393
rect 533674 78452 533738 80331
rect 534056 78452 534128 80331
rect 533674 41995 534128 78452
rect 535535 59924 535855 82391
rect 545937 84316 546950 84418
rect 545937 83115 546006 84316
rect 545937 82338 545974 83115
rect 546899 82515 546950 84316
rect 546865 82338 546950 82515
rect 552681 84259 553924 88193
rect 552681 82521 552784 84259
rect 553776 82521 553924 84259
rect 552681 82394 553924 82521
rect 545937 82265 546950 82338
rect 554170 81554 555098 89107
rect 552170 80626 555098 81554
rect 556570 84330 557114 84401
rect 556570 82460 556629 84330
rect 557062 82460 557114 84330
rect 566612 83547 567558 83651
rect 566612 83208 566647 83547
rect 567525 83208 567558 83547
rect 535535 58682 535562 59924
rect 535808 58682 535855 59924
rect 535535 58641 535855 58682
rect 536449 80392 536769 80396
rect 536449 80320 536936 80392
rect 536449 78457 536519 80320
rect 536865 78457 536936 80320
rect 552170 80271 553098 80626
rect 543134 80189 544731 80250
rect 543134 79844 543189 80189
rect 544669 79844 544731 80189
rect 543134 79804 543472 79844
rect 536449 78393 536936 78457
rect 536449 59928 536769 78393
rect 537339 75697 537482 79496
rect 543388 78615 543472 79804
rect 544433 79804 544731 79844
rect 544433 78615 544500 79804
rect 543388 78532 544500 78615
rect 552170 78565 552287 80271
rect 552970 78565 553098 80271
rect 552170 78405 553098 78565
rect 553970 80313 554514 80361
rect 553970 78446 554026 80313
rect 554459 78446 554514 80313
rect 538745 74308 539199 74386
rect 538745 69457 538810 74308
rect 539135 69457 539199 74308
rect 536449 58686 536487 59928
rect 536733 58686 536769 59928
rect 536449 58635 536769 58686
rect 537488 67322 537942 67408
rect 537488 62471 537554 67322
rect 537879 62471 537942 67322
rect 537488 57334 537942 62471
rect 533674 41736 533708 41995
rect 534074 41736 534128 41995
rect 533674 28437 534128 41736
rect 533674 28161 533717 28437
rect 534113 28161 534128 28437
rect 533674 21172 534128 28161
rect 536065 56880 537942 57334
rect 536065 35123 536519 56880
rect 538745 56249 539199 69457
rect 539719 67296 540744 76051
rect 539719 62457 539787 67296
rect 540637 62457 540744 67296
rect 539719 62094 540744 62457
rect 536065 34797 536094 35123
rect 536485 34797 536519 35123
rect 536065 21569 536519 34797
rect 536065 21250 536097 21569
rect 536489 21250 536519 21569
rect 536065 21111 536519 21250
rect 537306 55795 539199 56249
rect 537306 36166 537760 55795
rect 537306 35840 537333 36166
rect 537724 35840 537760 36166
rect 537306 22596 537760 35840
rect 537306 22277 537335 22596
rect 537727 22277 537760 22596
rect 537306 21141 537760 22277
rect 540307 17496 540572 47888
rect 540875 17863 541140 47888
rect 542038 33590 542166 73755
rect 542294 33167 542422 73235
rect 542550 33888 542678 72732
rect 553970 72555 554514 78446
rect 542806 34225 542934 72216
rect 551957 72011 554514 72555
rect 543062 46982 543190 68633
rect 543318 46718 543446 68130
rect 543574 47286 543702 67621
rect 543830 47521 543958 67133
rect 544086 60180 544214 66594
rect 544342 59829 544470 66077
rect 551957 55050 552501 72011
rect 556570 71158 557114 82460
rect 562850 82526 563986 82560
rect 562850 82178 562875 82526
rect 563960 82178 563986 82526
rect 551957 54794 551991 55050
rect 552467 54794 552501 55050
rect 551957 41808 552501 54794
rect 551957 41575 552005 41808
rect 552430 41575 552501 41808
rect 551957 28406 552501 41575
rect 551957 28194 551998 28406
rect 552437 28194 552501 28406
rect 551957 21111 552501 28194
rect 553198 70614 557114 71158
rect 557383 74307 557927 74399
rect 553198 54132 553742 70614
rect 557383 69934 557464 74307
rect 553198 53876 553227 54132
rect 553703 53876 553742 54132
rect 553198 40876 553742 53876
rect 553198 40643 553252 40876
rect 553677 40643 553742 40876
rect 553198 27515 553742 40643
rect 553198 27275 553259 27515
rect 553698 27275 553742 27515
rect 553198 21081 553742 27275
rect 556014 69463 557464 69934
rect 557847 69463 557927 74307
rect 556014 69390 557927 69463
rect 556014 49239 556558 69390
rect 558363 67325 558907 67394
rect 558363 62481 558449 67325
rect 558832 62481 558907 67325
rect 558363 62177 558907 62481
rect 556014 48910 556070 49239
rect 556495 48910 556558 49239
rect 556014 35981 556558 48910
rect 556014 35680 556063 35981
rect 556515 35680 556558 35981
rect 556014 22600 556558 35680
rect 556014 22285 556049 22600
rect 556515 22285 556558 22600
rect 556014 21050 556558 22285
rect 557285 61633 558907 62177
rect 562850 67301 563986 82178
rect 562850 62472 562936 67301
rect 563908 62472 563986 67301
rect 557285 48197 557829 61633
rect 562850 60715 563986 62472
rect 566612 74315 567558 83208
rect 566612 69459 566684 74315
rect 567369 69459 567558 74315
rect 562697 60665 564300 60715
rect 562697 60236 562759 60665
rect 564261 60236 564300 60665
rect 562697 60167 564300 60236
rect 557285 47868 557345 48197
rect 557770 47868 557829 48197
rect 557285 34932 557829 47868
rect 557285 34631 557338 34932
rect 557790 34631 557829 34932
rect 557285 21592 557829 34631
rect 557285 21277 557324 21592
rect 557790 21277 557829 21592
rect 546844 5674 547192 20228
rect 554920 6316 555294 20214
rect 518727 774 518780 2210
rect 519880 774 519927 2210
rect 557285 3138 557829 21277
rect 563199 9637 563388 17682
rect 563566 9985 563768 18042
rect 564256 10470 564556 21524
rect 564856 10879 565156 20404
rect 565456 11288 565756 61110
rect 566056 11804 566356 60044
rect 566612 59030 567558 69459
rect 566612 58523 566623 59030
rect 567534 58523 567558 59030
rect 566612 58467 567558 58523
rect 570962 67340 571354 75526
rect 570962 66204 571006 67340
rect 571316 66204 571354 67340
rect 566656 12354 566956 48710
rect 567256 12727 567556 51914
rect 567856 13154 568156 46872
rect 568456 13582 568756 44556
rect 569056 14068 569356 35442
rect 569656 14442 569956 34798
rect 570256 14957 570556 33530
rect 570962 33212 571354 66204
rect 570856 15377 571156 28008
rect 571856 15794 572156 80744
rect 572456 34178 572756 81739
rect 573056 55816 573356 94580
rect 573656 94288 573665 95095
rect 573719 94288 573956 95095
rect 573656 76164 573956 94288
rect 570856 15249 572272 15377
rect 570256 14829 571760 14957
rect 569656 14314 571248 14442
rect 569056 13940 570736 14068
rect 568456 13454 570224 13582
rect 567856 13026 569712 13154
rect 567256 12599 569200 12727
rect 566656 12226 568688 12354
rect 566056 11676 567664 11804
rect 565456 11160 567152 11288
rect 564856 10751 566640 10879
rect 564256 10342 566128 10470
rect 563566 9857 565616 9985
rect 563199 9509 565104 9637
rect 562016 3941 562144 8461
rect 562528 4306 562656 8968
rect 563040 4671 563168 8559
rect 563552 5125 563680 8160
rect 564064 5598 564192 7761
rect 564064 5470 564592 5598
rect 563552 4997 564080 5125
rect 563040 4543 563568 4671
rect 562528 4178 563056 4306
rect 562016 3813 562544 3941
rect 557285 2170 557330 3138
rect 557790 2170 557829 3138
rect 557285 2132 557829 2170
rect 518727 640 519927 774
rect 562156 0 562284 3179
rect 562416 0 562544 3813
rect 562668 0 562796 3179
rect 562928 0 563056 4178
rect 563180 0 563308 3179
rect 563440 0 563568 4543
rect 563692 0 563820 3179
rect 563952 0 564080 4997
rect 564204 0 564332 3179
rect 564464 0 564592 5470
rect 564716 0 564844 3179
rect 564976 0 565104 9509
rect 565228 0 565356 3179
rect 565488 0 565616 9857
rect 565740 0 565868 3179
rect 566000 0 566128 10342
rect 566260 0 566388 3179
rect 566512 0 566640 10751
rect 566772 0 566900 3179
rect 567024 0 567152 11160
rect 567284 0 567412 3179
rect 567536 0 567664 11676
rect 567796 0 567924 3179
rect 568048 0 568176 9580
rect 568308 0 568436 3179
rect 568560 0 568688 12226
rect 568820 0 568948 3179
rect 569072 0 569200 12599
rect 569332 0 569460 3179
rect 569584 0 569712 13026
rect 569844 0 569972 3179
rect 570096 0 570224 13454
rect 570356 0 570484 3179
rect 570608 0 570736 13940
rect 570868 0 570996 3179
rect 571120 0 571248 14314
rect 571380 0 571508 3179
rect 571632 0 571760 14829
rect 571892 0 572020 3179
rect 572144 0 572272 15249
rect 572676 12214 573010 33536
rect 572404 0 572532 3179
<< rmetal4 >>
rect 354960 3068 355088 3114
rect 355472 3068 355600 3114
rect 355984 3068 356112 3114
rect 356496 3068 356624 3114
rect 357008 3068 357136 3114
rect 357520 3068 357648 3114
rect 358032 3068 358160 3114
rect 358544 3068 358672 3114
rect 359056 3068 359184 3114
rect 359568 3068 359696 3114
rect 360080 3068 360208 3114
rect 360592 3068 360720 3114
rect 361104 3068 361232 3114
rect 361616 3068 361744 3114
rect 362128 3068 362256 3114
rect 362640 3068 362768 3114
<< via4 >>
rect 25090 83562 25749 84356
rect 25090 83300 25531 83562
rect 25531 83300 25749 83562
rect 25090 82430 25749 83300
rect 15421 69442 16093 74356
rect 11043 64365 14614 65195
rect 20258 62506 20918 67331
rect 29921 78434 30580 80360
rect 37821 82462 38379 84315
rect 37010 69435 37641 74322
rect 38721 78461 39238 80323
rect 39559 62500 40217 67339
rect 40801 69472 41224 74319
rect 43708 69482 44464 74274
rect 46784 82470 47234 84312
rect 41507 62466 42011 67339
rect 46174 78464 46624 80306
rect 45004 62518 45760 67310
rect 83914 69498 84573 74312
rect 91979 69425 92280 74308
rect 83875 58740 84621 61116
rect 81321 11629 82276 13072
rect 85099 62454 85769 67220
rect 90989 62474 91290 67357
rect 96440 82461 96740 84319
rect 97352 78446 97652 80304
rect 131380 110345 132311 111807
rect 118373 69535 120308 74180
rect 130258 82434 130778 84334
rect 129052 78442 129572 80342
rect 127814 69488 128339 74293
rect 121918 62593 123526 67196
rect 126488 62493 127013 67298
rect 132983 107951 133914 109413
rect 139578 82437 140216 84335
rect 140461 80003 141130 80339
rect 140461 79863 141130 80003
rect 140461 78428 141130 79863
rect 141534 69463 142314 74335
rect 155647 82449 156028 84353
rect 154843 78438 155224 80342
rect 153620 69472 155025 74319
rect 142726 62453 143472 67337
rect 150178 62514 151580 67300
rect 161026 82456 161275 84342
rect 182529 82473 183204 84328
rect 160495 78449 160744 80335
rect 159333 69523 159746 74294
rect 160173 62500 160653 67284
rect 82751 8021 83706 9464
rect 91118 3174 91406 4643
rect 123625 3181 123912 4661
rect 90590 765 90878 2234
rect 193333 82436 193619 84330
rect 184167 78472 185074 80307
rect 186750 78451 187269 80328
rect 193869 78449 194155 80343
rect 191297 69495 191872 74303
rect 189982 62495 190557 67303
rect 195491 69507 195955 74320
rect 199850 82511 200371 84345
rect 198882 80135 199386 80358
rect 198882 79994 199386 80135
rect 198882 78457 199386 79994
rect 203025 82447 203443 84336
rect 194459 62511 194939 67249
rect 212614 69514 213958 74261
rect 207583 62469 208056 67295
rect 209202 62505 210546 67252
rect 230551 69592 232344 74231
rect 132718 8142 133480 9650
rect 131510 5738 132272 7246
rect 124153 757 124440 2237
rect 156181 3258 157163 4622
rect 148608 819 149590 2183
rect 172217 759 172892 2245
rect 173431 3176 174106 4662
rect 247420 69468 248462 74305
rect 234444 62540 238960 67234
rect 245474 62489 246432 67297
rect 215109 3227 216072 4611
rect 207569 807 208532 2191
rect 230517 759 231189 2250
rect 253359 69491 256333 74267
rect 249437 62494 252411 67270
rect 257364 69460 257711 74319
rect 268502 82442 268889 84351
rect 258542 62522 262334 67274
rect 267689 69489 267990 74348
rect 266840 62501 267165 67328
rect 272385 82464 272639 84347
rect 273026 78456 273529 80334
rect 277546 69450 277912 74336
rect 275169 62522 275693 67273
rect 279860 69470 280452 74306
rect 282083 62444 282449 67330
rect 231731 3176 232396 4664
rect 254124 3198 254704 4660
rect 277360 3262 278170 4628
rect 251034 751 251979 2235
rect 286644 82522 287651 84302
rect 298712 82446 299135 84349
rect 286652 3247 287645 4600
rect 288414 78505 289421 80285
rect 279768 786 280605 2213
rect 299757 78472 300134 80328
rect 290546 69512 291120 74305
rect 293782 69482 294150 74317
rect 311386 82474 312087 84307
rect 311397 75481 312080 77590
rect 303458 69526 308006 74274
rect 313130 69514 317694 74234
rect 292652 62487 293020 67322
rect 320991 82442 321227 84344
rect 321887 78667 322125 80353
rect 445406 110390 449996 111737
rect 450659 108010 455028 109358
rect 319884 69448 320146 74324
rect 346037 69476 346312 74285
rect 319016 62470 319300 67334
rect 345399 62459 345859 67319
rect 290503 59454 291181 61397
rect 346554 62455 346815 67296
rect 352700 69569 353645 74295
rect 352418 62486 353986 67250
rect 347668 50652 351477 53453
rect 288423 820 289416 2173
rect 339670 14892 340952 15312
rect 339692 11465 340974 11885
rect 338746 3172 339105 4669
rect 341501 3176 341760 4673
rect 294538 796 294988 2206
rect 341930 747 342210 2237
rect 366319 82451 366642 84329
rect 363842 62496 364730 67288
rect 365384 78476 365659 80321
rect 365904 78432 366152 80311
rect 367001 82450 367267 84346
rect 371627 82450 371893 84346
rect 370530 78432 370778 80311
rect 374726 82435 375181 84318
rect 376253 82450 376519 84346
rect 375516 80126 376086 80350
rect 375516 79999 376086 80126
rect 375516 78432 376086 79999
rect 368232 69414 368531 74363
rect 380879 82450 381145 84346
rect 372858 69414 373157 74363
rect 369876 62448 370126 67349
rect 372355 62506 373406 67295
rect 374411 69477 375214 74290
rect 376090 69459 376822 74328
rect 377484 69414 377783 74363
rect 378163 62448 378932 67323
rect 363198 20548 363516 21284
rect 379982 78432 380230 80311
rect 385474 82438 386053 84350
rect 384408 78432 385036 80337
rect 382110 69414 382409 74363
rect 379128 62448 379378 67349
rect 383754 62448 384004 67349
rect 382998 50614 383893 53463
rect 364589 15024 365295 16947
rect 368294 44750 369665 45515
rect 388948 82465 389318 84328
rect 389034 78432 389282 80311
rect 389905 78524 390347 80315
rect 386736 69414 387035 74363
rect 388380 62448 388630 67349
rect 384400 39126 385734 39680
rect 391692 69422 391938 74343
rect 395377 82442 395670 84285
rect 399383 82450 399649 84346
rect 393607 78434 393862 78889
rect 394948 78459 395252 80338
rect 396692 78431 397253 80346
rect 393729 69498 394202 74321
rect 393277 62461 393531 67327
rect 395988 69414 396287 74363
rect 394738 62485 395227 67323
rect 398286 78432 398534 80311
rect 403823 82436 404281 84347
rect 402912 78432 403367 80341
rect 400614 69414 400913 74363
rect 397632 62448 397882 67349
rect 402258 62448 402508 67349
rect 408635 82450 408901 84346
rect 407538 78432 407786 80311
rect 413261 82450 413527 84346
rect 412164 78432 412412 80311
rect 417887 82450 418153 84346
rect 416790 78432 417038 80311
rect 422513 82450 422779 84346
rect 421416 78432 421664 80311
rect 424351 82430 424599 84339
rect 405240 69414 405539 74363
rect 409866 69414 410165 74363
rect 406884 62448 407134 67349
rect 414492 69414 414791 74363
rect 411510 62448 411760 67349
rect 419118 69414 419417 74363
rect 416136 62448 416386 67349
rect 422587 69456 423195 74339
rect 420762 62448 421012 67349
rect 421550 62471 422153 67324
rect 414932 60678 415612 61829
rect 389744 50582 390995 53468
rect 391494 45614 392733 48413
rect 423744 69414 424043 74363
rect 427404 82476 427681 84189
rect 424822 78438 425070 80347
rect 426042 78432 426290 80311
rect 427942 78463 428243 80342
rect 431765 82450 432031 84346
rect 427997 69455 428235 74338
rect 425388 62448 425638 67349
rect 430968 78432 431216 80311
rect 429574 69452 430005 74290
rect 428531 62479 429041 67316
rect 435287 82453 435737 84337
rect 436391 82450 436657 84346
rect 434297 78449 434747 80333
rect 435294 78432 435542 80311
rect 441017 82450 441283 84346
rect 440090 78432 440338 80311
rect 445643 82450 445909 84346
rect 444716 78432 444964 80311
rect 450269 82450 450535 84346
rect 449172 78432 449420 80311
rect 451692 82445 452265 84338
rect 450780 80303 451361 80358
rect 450780 80161 451361 80303
rect 450780 78430 451361 80161
rect 434031 70845 434276 74329
rect 430327 62443 430568 67349
rect 405504 45583 406457 48473
rect 431483 62472 432140 67324
rect 437622 69414 437921 74363
rect 435109 62462 435349 67346
rect 442248 69414 442547 74363
rect 439266 62448 439516 67349
rect 446874 69414 447173 74363
rect 443892 62448 444142 67349
rect 451500 69414 451799 74363
rect 448518 62448 448768 67349
rect 454895 82450 455161 84346
rect 453968 78432 454216 80311
rect 459521 82450 459787 84346
rect 458624 78432 458872 80311
rect 464147 82450 464413 84346
rect 463150 78432 463398 80311
rect 456126 69414 456425 74363
rect 453044 62448 453294 67349
rect 460752 69414 461051 74363
rect 457770 62448 458020 67349
rect 464711 69463 464949 74342
rect 462196 62448 462446 67349
rect 486280 86228 490240 89522
rect 468773 82450 469039 84346
rect 467876 78432 468124 80311
rect 473399 82450 473665 84346
rect 472502 78432 472750 80311
rect 470004 69414 470303 74363
rect 465312 62510 467131 67277
rect 478025 84345 478291 84346
rect 478025 82450 478720 84345
rect 476801 78423 477563 80342
rect 474098 69572 475813 74237
rect 471248 62448 471498 67349
rect 476174 62448 476424 67349
rect 482651 82450 482917 84346
rect 481754 78432 482002 80311
rect 479256 69414 479555 74363
rect 487277 82450 487543 84346
rect 486380 78432 486628 80311
rect 480900 62448 481150 67349
rect 484043 69527 485525 74249
rect 491006 78432 491254 80311
rect 491903 82450 492169 84346
rect 496529 82450 496795 84346
rect 495632 78432 495880 80311
rect 499199 82442 499453 84323
rect 498269 78443 498514 80325
rect 499958 78432 500206 80311
rect 501155 83150 501421 84346
rect 501155 82450 501407 83150
rect 501407 82450 501421 83150
rect 488817 69518 490270 74302
rect 486318 62481 486562 67310
rect 487006 62510 488459 67294
rect 493134 69414 493433 74363
rect 490841 62471 491077 67346
rect 494578 62448 494828 67349
rect 496534 69510 497987 74294
rect 498357 62507 499810 67291
rect 502386 69414 502685 74363
rect 500401 62445 500662 67353
rect 507329 69529 508782 74313
rect 503780 62448 504030 67349
rect 505496 62478 506949 67262
rect 511154 85727 515114 89021
rect 532883 82455 533201 83634
rect 515008 69510 516461 74294
rect 509143 62497 510596 67281
rect 516863 62497 518316 67281
rect 530609 69458 530860 74316
rect 529618 62466 529869 67324
rect 521477 45689 525395 48410
rect 475586 18455 478387 19501
rect 479182 18553 480378 20475
rect 365875 15047 366581 16970
rect 363655 13435 364110 14724
rect 364566 11594 365310 13158
rect 365865 9755 366609 11319
rect 487572 10414 488240 10794
rect 475597 6385 476706 7697
rect 364588 770 365003 2226
rect 475597 824 476706 2136
rect 490718 3276 491898 4624
rect 494902 3202 496002 4638
rect 485221 843 486580 2202
rect 500288 774 501388 2210
rect 509316 3217 510361 4588
rect 513408 3198 514508 4634
rect 503942 801 504987 2172
rect 535463 82458 535798 84314
rect 533738 78452 534056 80331
rect 546006 83115 546899 84316
rect 546006 82515 546865 83115
rect 546865 82515 546899 83115
rect 552784 82521 553776 84259
rect 556629 82460 557062 84330
rect 536519 78457 536865 80320
rect 543472 79844 544433 80189
rect 543472 78615 544433 79844
rect 552287 78565 552970 80271
rect 554026 78446 554459 80313
rect 538810 69457 539135 74308
rect 537554 62471 537879 67322
rect 539787 62457 540637 67296
rect 557464 69463 557847 74307
rect 558449 62481 558832 67325
rect 562936 62472 563908 67301
rect 566684 69459 567369 74315
rect 518780 774 519880 2210
rect 571006 66204 571316 67340
<< metal5 >>
rect 131284 111807 450217 111876
rect 131284 110345 131380 111807
rect 132311 111737 450217 111807
rect 132311 110390 445406 111737
rect 449996 110390 450217 111737
rect 132311 110345 450217 110390
rect 131284 110276 450217 110345
rect -4 109022 6832 110022
rect 132876 109413 455228 109476
rect -4 107022 19277 109022
rect 132876 107951 132983 109413
rect 133914 109358 455228 109413
rect 133914 108010 450659 109358
rect 455028 108010 455228 109358
rect 563080 109169 574622 110022
rect 133914 107951 455228 108010
rect 132876 107876 455228 107951
rect -4 103022 14337 105022
rect -4 102022 6832 103022
rect 349 93220 7988 93540
rect 0 92220 5620 92540
rect 12337 80390 14337 103022
rect 17277 84390 19277 107022
rect 558232 107024 574622 109169
rect 486148 89522 501016 89656
rect 486148 86228 486280 89522
rect 490240 89156 501016 89522
rect 490240 89021 515268 89156
rect 490240 86228 511154 89021
rect 486148 86098 511154 86228
rect 496961 85727 511154 86098
rect 515114 85727 515268 89021
rect 496961 85598 515268 85727
rect 558232 84390 560232 107024
rect 563080 107022 574622 107024
rect 17277 84356 560232 84390
rect 17277 82430 25090 84356
rect 25749 84353 560232 84356
rect 25749 84335 155647 84353
rect 25749 84334 139578 84335
rect 25749 84319 130258 84334
rect 25749 84315 96440 84319
rect 25749 82462 37821 84315
rect 38379 84312 96440 84315
rect 38379 82470 46784 84312
rect 47234 82470 96440 84312
rect 38379 82462 96440 82470
rect 25749 82461 96440 82462
rect 96740 82461 130258 84319
rect 25749 82434 130258 82461
rect 130778 82437 139578 84334
rect 140216 82449 155647 84335
rect 156028 84351 560232 84353
rect 156028 84345 268502 84351
rect 156028 84342 199850 84345
rect 156028 82456 161026 84342
rect 161275 84330 199850 84342
rect 161275 84328 193333 84330
rect 161275 82473 182529 84328
rect 183204 82473 193333 84328
rect 161275 82456 193333 82473
rect 156028 82449 193333 82456
rect 140216 82437 193333 82449
rect 130778 82436 193333 82437
rect 193619 82511 199850 84330
rect 200371 84336 268502 84345
rect 200371 82511 203025 84336
rect 193619 82447 203025 82511
rect 203443 82447 268502 84336
rect 193619 82442 268502 82447
rect 268889 84350 560232 84351
rect 268889 84349 385474 84350
rect 268889 84347 298712 84349
rect 268889 82464 272385 84347
rect 272639 84302 298712 84347
rect 272639 82522 286644 84302
rect 287651 82522 298712 84302
rect 272639 82464 298712 82522
rect 268889 82446 298712 82464
rect 299135 84346 385474 84349
rect 299135 84344 367001 84346
rect 299135 84307 320991 84344
rect 299135 82474 311386 84307
rect 312087 82474 320991 84307
rect 299135 82446 320991 82474
rect 268889 82442 320991 82446
rect 321227 84329 367001 84344
rect 321227 82451 366319 84329
rect 366642 82451 367001 84329
rect 321227 82450 367001 82451
rect 367267 82450 371627 84346
rect 371893 84318 376253 84346
rect 371893 82450 374726 84318
rect 321227 82442 374726 82450
rect 193619 82436 374726 82442
rect 130778 82435 374726 82436
rect 375181 82450 376253 84318
rect 376519 82450 380879 84346
rect 381145 82450 385474 84346
rect 375181 82438 385474 82450
rect 386053 84347 560232 84350
rect 386053 84346 403823 84347
rect 386053 84328 399383 84346
rect 386053 82465 388948 84328
rect 389318 84285 399383 84328
rect 389318 82465 395377 84285
rect 386053 82442 395377 82465
rect 395670 82450 399383 84285
rect 399649 82450 403823 84346
rect 395670 82442 403823 82450
rect 386053 82438 403823 82442
rect 375181 82436 403823 82438
rect 404281 84346 560232 84347
rect 404281 82450 408635 84346
rect 408901 82450 413261 84346
rect 413527 82450 417887 84346
rect 418153 82450 422513 84346
rect 422779 84339 431765 84346
rect 422779 82450 424351 84339
rect 404281 82436 424351 82450
rect 375181 82435 424351 82436
rect 130778 82434 424351 82435
rect 25749 82430 424351 82434
rect 424599 84189 431765 84339
rect 424599 82476 427404 84189
rect 427681 82476 431765 84189
rect 424599 82450 431765 82476
rect 432031 84337 436391 84346
rect 432031 82453 435287 84337
rect 435737 82453 436391 84337
rect 432031 82450 436391 82453
rect 436657 82450 441017 84346
rect 441283 82450 445643 84346
rect 445909 82450 450269 84346
rect 450535 84338 454895 84346
rect 450535 82450 451692 84338
rect 424599 82445 451692 82450
rect 452265 82450 454895 84338
rect 455161 82450 459521 84346
rect 459787 82450 464147 84346
rect 464413 82450 468773 84346
rect 469039 82450 473399 84346
rect 473665 82450 478025 84346
rect 478291 84345 482651 84346
rect 478720 82450 482651 84345
rect 482917 82450 487277 84346
rect 487543 82450 491903 84346
rect 492169 82450 496529 84346
rect 496795 84323 501155 84346
rect 496795 82450 499199 84323
rect 452265 82445 499199 82450
rect 424599 82442 499199 82445
rect 499453 82450 501155 84323
rect 501421 84330 560232 84346
rect 501421 84316 556629 84330
rect 501421 84314 546006 84316
rect 501421 83634 535463 84314
rect 501421 82455 532883 83634
rect 533201 82458 535463 83634
rect 535798 82515 546006 84314
rect 546899 84259 556629 84316
rect 546899 82521 552784 84259
rect 553776 82521 556629 84259
rect 546899 82515 556629 82521
rect 535798 82460 556629 82515
rect 557062 82460 560232 84330
rect 535798 82458 560232 82460
rect 533201 82455 560232 82458
rect 501421 82450 560232 82455
rect 499453 82442 560232 82450
rect 424599 82430 560232 82442
rect 17277 82390 560232 82430
rect 561798 105022 563128 105023
rect 561798 102022 574622 105022
rect 561798 80390 563798 102022
rect 12337 80360 563798 80390
rect 12337 78434 29921 80360
rect 30580 80358 563798 80360
rect 30580 80343 198882 80358
rect 30580 80342 193869 80343
rect 30580 80323 129052 80342
rect 30580 78461 38721 80323
rect 39238 80306 129052 80323
rect 39238 78464 46174 80306
rect 46624 80304 129052 80306
rect 46624 78464 97352 80304
rect 39238 78461 97352 78464
rect 30580 78446 97352 78461
rect 97652 78446 129052 80304
rect 30580 78442 129052 78446
rect 129572 80339 154843 80342
rect 129572 78442 140461 80339
rect 30580 78434 140461 78442
rect 12337 78428 140461 78434
rect 141130 78438 154843 80339
rect 155224 80335 193869 80342
rect 155224 78449 160495 80335
rect 160744 80328 193869 80335
rect 160744 80307 186750 80328
rect 160744 78472 184167 80307
rect 185074 78472 186750 80307
rect 160744 78451 186750 78472
rect 187269 78451 193869 80328
rect 160744 78449 193869 78451
rect 194155 78457 198882 80343
rect 199386 80353 450780 80358
rect 199386 80334 321887 80353
rect 199386 78457 273026 80334
rect 194155 78456 273026 78457
rect 273529 80328 321887 80334
rect 273529 80285 299757 80328
rect 273529 78505 288414 80285
rect 289421 78505 299757 80285
rect 273529 78472 299757 78505
rect 300134 78667 321887 80328
rect 322125 80350 450780 80353
rect 322125 80321 375516 80350
rect 322125 78667 365384 80321
rect 300134 78476 365384 78667
rect 365659 80311 375516 80321
rect 365659 78476 365904 80311
rect 300134 78472 365904 78476
rect 273529 78456 365904 78472
rect 194155 78449 365904 78456
rect 155224 78438 365904 78449
rect 141130 78432 365904 78438
rect 366152 78432 370530 80311
rect 370778 78432 375516 80311
rect 376086 80347 450780 80350
rect 376086 80346 424822 80347
rect 376086 80338 396692 80346
rect 376086 80337 394948 80338
rect 376086 80311 384408 80337
rect 376086 78432 379982 80311
rect 380230 78432 384408 80311
rect 385036 80315 394948 80337
rect 385036 80311 389905 80315
rect 385036 78432 389034 80311
rect 389282 78524 389905 80311
rect 390347 78889 394948 80315
rect 390347 78524 393607 78889
rect 389282 78434 393607 78524
rect 393862 78459 394948 78889
rect 395252 78459 396692 80338
rect 393862 78434 396692 78459
rect 389282 78432 396692 78434
rect 141130 78431 396692 78432
rect 397253 80341 424822 80346
rect 397253 80311 402912 80341
rect 397253 78432 398286 80311
rect 398534 78432 402912 80311
rect 403367 80311 424822 80341
rect 403367 78432 407538 80311
rect 407786 78432 412164 80311
rect 412412 78432 416790 80311
rect 417038 78432 421416 80311
rect 421664 78438 424822 80311
rect 425070 80342 450780 80347
rect 425070 80311 427942 80342
rect 425070 78438 426042 80311
rect 421664 78432 426042 78438
rect 426290 78463 427942 80311
rect 428243 80333 450780 80342
rect 428243 80311 434297 80333
rect 428243 78463 430968 80311
rect 426290 78432 430968 78463
rect 431216 78449 434297 80311
rect 434747 80311 450780 80333
rect 434747 78449 435294 80311
rect 431216 78432 435294 78449
rect 435542 78432 440090 80311
rect 440338 78432 444716 80311
rect 444964 78432 449172 80311
rect 449420 78432 450780 80311
rect 397253 78431 450780 78432
rect 141130 78430 450780 78431
rect 451361 80342 563798 80358
rect 451361 80311 476801 80342
rect 451361 78432 453968 80311
rect 454216 78432 458624 80311
rect 458872 78432 463150 80311
rect 463398 78432 467876 80311
rect 468124 78432 472502 80311
rect 472750 78432 476801 80311
rect 451361 78430 476801 78432
rect 141130 78428 476801 78430
rect 12337 78423 476801 78428
rect 477563 80331 563798 80342
rect 477563 80325 533738 80331
rect 477563 80311 498269 80325
rect 477563 78432 481754 80311
rect 482002 78432 486380 80311
rect 486628 78432 491006 80311
rect 491254 78432 495632 80311
rect 495880 78443 498269 80311
rect 498514 80311 533738 80325
rect 498514 78443 499958 80311
rect 495880 78432 499958 78443
rect 500206 78452 533738 80311
rect 534056 80320 563798 80331
rect 534056 78457 536519 80320
rect 536865 80313 563798 80320
rect 536865 80271 554026 80313
rect 536865 80189 552287 80271
rect 536865 78615 543472 80189
rect 544433 78615 552287 80189
rect 536865 78565 552287 78615
rect 552970 78565 554026 80271
rect 536865 78457 554026 78565
rect 534056 78452 554026 78457
rect 500206 78446 554026 78452
rect 554459 78446 563798 80313
rect 500206 78432 563798 78446
rect 477563 78423 563798 78432
rect 12337 78390 563798 78423
rect 311310 77590 312178 77702
rect 311310 75481 311397 77590
rect 312080 77092 312178 77590
rect 312080 76675 345371 77092
rect 312080 75481 312178 76675
rect 573641 76200 574620 76520
rect 311310 75373 312178 75481
rect 570949 75198 574276 75518
rect 10930 74363 567508 74390
rect 10930 74356 368232 74363
rect 349 72220 7990 72540
rect 0 71220 5620 71540
rect 10930 69442 15421 74356
rect 16093 74348 368232 74356
rect 16093 74335 267689 74348
rect 16093 74322 141534 74335
rect 16093 69442 37010 74322
rect 10930 69435 37010 69442
rect 37641 74319 141534 74322
rect 37641 69472 40801 74319
rect 41224 74312 141534 74319
rect 41224 74274 83914 74312
rect 41224 69482 43708 74274
rect 44464 69498 83914 74274
rect 84573 74308 141534 74312
rect 84573 69498 91979 74308
rect 44464 69482 91979 69498
rect 41224 69472 91979 69482
rect 37641 69435 91979 69472
rect 10930 69425 91979 69435
rect 92280 74293 141534 74308
rect 92280 74180 127814 74293
rect 92280 69535 118373 74180
rect 120308 69535 127814 74180
rect 92280 69488 127814 69535
rect 128339 69488 141534 74293
rect 92280 69463 141534 69488
rect 142314 74320 267689 74335
rect 142314 74319 195491 74320
rect 142314 69472 153620 74319
rect 155025 74303 195491 74319
rect 155025 74294 191297 74303
rect 155025 69523 159333 74294
rect 159746 69523 191297 74294
rect 155025 69495 191297 69523
rect 191872 69507 195491 74303
rect 195955 74319 267689 74320
rect 195955 74305 257364 74319
rect 195955 74261 247420 74305
rect 195955 69514 212614 74261
rect 213958 74231 247420 74261
rect 213958 69592 230551 74231
rect 232344 69592 247420 74231
rect 213958 69514 247420 69592
rect 195955 69507 247420 69514
rect 191872 69495 247420 69507
rect 155025 69472 247420 69495
rect 142314 69468 247420 69472
rect 248462 74267 257364 74305
rect 248462 69491 253359 74267
rect 256333 69491 257364 74267
rect 248462 69468 257364 69491
rect 142314 69463 257364 69468
rect 92280 69460 257364 69463
rect 257711 69489 267689 74319
rect 267990 74336 368232 74348
rect 267990 69489 277546 74336
rect 257711 69460 277546 69489
rect 92280 69450 277546 69460
rect 277912 74324 368232 74336
rect 277912 74317 319884 74324
rect 277912 74306 293782 74317
rect 277912 69470 279860 74306
rect 280452 74305 293782 74306
rect 280452 69512 290546 74305
rect 291120 69512 293782 74305
rect 280452 69482 293782 69512
rect 294150 74274 319884 74317
rect 294150 69526 303458 74274
rect 308006 74234 319884 74274
rect 308006 69526 313130 74234
rect 294150 69514 313130 69526
rect 317694 69514 319884 74234
rect 294150 69482 319884 69514
rect 280452 69470 319884 69482
rect 277912 69450 319884 69470
rect 92280 69448 319884 69450
rect 320146 74295 368232 74324
rect 320146 74285 352700 74295
rect 320146 69476 346037 74285
rect 346312 69569 352700 74285
rect 353645 69569 368232 74295
rect 346312 69476 368232 69569
rect 320146 69448 368232 69476
rect 92280 69425 368232 69448
rect 10930 69414 368232 69425
rect 368531 69414 372858 74363
rect 373157 74328 377484 74363
rect 373157 74290 376090 74328
rect 373157 69477 374411 74290
rect 375214 69477 376090 74290
rect 373157 69459 376090 69477
rect 376822 69459 377484 74328
rect 373157 69414 377484 69459
rect 377783 69414 382110 74363
rect 382409 69414 386736 74363
rect 387035 74343 395988 74363
rect 387035 69422 391692 74343
rect 391938 74321 395988 74343
rect 391938 69498 393729 74321
rect 394202 69498 395988 74321
rect 391938 69422 395988 69498
rect 387035 69414 395988 69422
rect 396287 69414 400614 74363
rect 400913 69414 405240 74363
rect 405539 69414 409866 74363
rect 410165 69414 414492 74363
rect 414791 69414 419118 74363
rect 419417 74339 423744 74363
rect 419417 69456 422587 74339
rect 423195 69456 423744 74339
rect 419417 69414 423744 69456
rect 424043 74338 437622 74363
rect 424043 69455 427997 74338
rect 428235 74329 437622 74338
rect 428235 74290 434031 74329
rect 428235 69455 429574 74290
rect 424043 69452 429574 69455
rect 430005 70845 434031 74290
rect 434276 70845 437622 74329
rect 430005 69452 437622 70845
rect 424043 69414 437622 69452
rect 437921 69414 442248 74363
rect 442547 69414 446874 74363
rect 447173 69414 451500 74363
rect 451799 69414 456126 74363
rect 456425 69414 460752 74363
rect 461051 74342 470004 74363
rect 461051 69463 464711 74342
rect 464949 69463 470004 74342
rect 461051 69414 470004 69463
rect 470303 74237 479256 74363
rect 470303 69572 474098 74237
rect 475813 69572 479256 74237
rect 470303 69414 479256 69572
rect 479555 74302 493134 74363
rect 479555 74249 488817 74302
rect 479555 69527 484043 74249
rect 485525 69527 488817 74249
rect 479555 69518 488817 69527
rect 490270 69518 493134 74302
rect 479555 69414 493134 69518
rect 493433 74294 502386 74363
rect 493433 69510 496534 74294
rect 497987 69510 502386 74294
rect 493433 69414 502386 69510
rect 502685 74316 567508 74363
rect 502685 74313 530609 74316
rect 502685 69529 507329 74313
rect 508782 74294 530609 74313
rect 508782 69529 515008 74294
rect 502685 69510 515008 69529
rect 516461 69510 530609 74294
rect 502685 69458 530609 69510
rect 530860 74315 567508 74316
rect 530860 74308 566684 74315
rect 530860 69458 538810 74308
rect 502685 69457 538810 69458
rect 539135 74307 566684 74308
rect 539135 69463 557464 74307
rect 557847 69463 566684 74307
rect 539135 69459 566684 69463
rect 567369 69459 567508 74315
rect 539135 69457 567508 69459
rect 502685 69414 567508 69457
rect 10930 69390 567508 69414
rect 298734 68934 299575 69390
rect 331910 68984 332631 69390
rect 293314 68373 318762 68934
rect 319614 68422 345148 68984
rect 10930 67357 571358 67390
rect 10930 67339 90989 67357
rect 10930 67331 39559 67339
rect 10930 65195 20258 67331
rect 10930 64365 11043 65195
rect 14614 64365 20258 65195
rect 10930 62506 20258 64365
rect 20918 62506 39559 67331
rect 10930 62500 39559 62506
rect 40217 62500 41507 67339
rect 10930 62466 41507 62500
rect 42011 67310 90989 67339
rect 42011 62518 45004 67310
rect 45760 67220 90989 67310
rect 45760 62518 85099 67220
rect 42011 62466 85099 62518
rect 10930 62454 85099 62466
rect 85769 62474 90989 67220
rect 91290 67353 571358 67357
rect 91290 67349 500401 67353
rect 91290 67337 369876 67349
rect 91290 67298 142726 67337
rect 91290 67196 126488 67298
rect 91290 62593 121918 67196
rect 123526 62593 126488 67196
rect 91290 62493 126488 62593
rect 127013 62493 142726 67298
rect 91290 62474 142726 62493
rect 85769 62454 142726 62474
rect 10930 62453 142726 62454
rect 143472 67334 369876 67337
rect 143472 67330 319016 67334
rect 143472 67328 282083 67330
rect 143472 67303 266840 67328
rect 143472 67300 189982 67303
rect 143472 62514 150178 67300
rect 151580 67284 189982 67300
rect 151580 62514 160173 67284
rect 143472 62500 160173 62514
rect 160653 62500 189982 67284
rect 143472 62495 189982 62500
rect 190557 67297 266840 67303
rect 190557 67295 245474 67297
rect 190557 67249 207583 67295
rect 190557 62511 194459 67249
rect 194939 62511 207583 67249
rect 190557 62495 207583 62511
rect 143472 62469 207583 62495
rect 208056 67252 245474 67295
rect 208056 62505 209202 67252
rect 210546 67234 245474 67252
rect 210546 62540 234444 67234
rect 238960 62540 245474 67234
rect 210546 62505 245474 62540
rect 208056 62489 245474 62505
rect 246432 67274 266840 67297
rect 246432 67270 258542 67274
rect 246432 62494 249437 67270
rect 252411 62522 258542 67270
rect 262334 62522 266840 67274
rect 252411 62501 266840 62522
rect 267165 67273 282083 67328
rect 267165 62522 275169 67273
rect 275693 62522 282083 67273
rect 267165 62501 282083 62522
rect 252411 62494 282083 62501
rect 246432 62489 282083 62494
rect 208056 62469 282083 62489
rect 143472 62453 282083 62469
rect 10930 62444 282083 62453
rect 282449 67322 319016 67330
rect 282449 62487 292652 67322
rect 293020 62487 319016 67322
rect 282449 62470 319016 62487
rect 319300 67319 369876 67334
rect 319300 62470 345399 67319
rect 282449 62459 345399 62470
rect 345859 67296 369876 67319
rect 345859 62459 346554 67296
rect 282449 62455 346554 62459
rect 346815 67288 369876 67296
rect 346815 67250 363842 67288
rect 346815 62486 352418 67250
rect 353986 62496 363842 67250
rect 364730 62496 369876 67288
rect 353986 62486 369876 62496
rect 346815 62455 369876 62486
rect 282449 62448 369876 62455
rect 370126 67323 379128 67349
rect 370126 67295 378163 67323
rect 370126 62506 372355 67295
rect 373406 62506 378163 67295
rect 370126 62448 378163 62506
rect 378932 62448 379128 67323
rect 379378 62448 383754 67349
rect 384004 62448 388380 67349
rect 388630 67327 397632 67349
rect 388630 62461 393277 67327
rect 393531 67323 397632 67327
rect 393531 62485 394738 67323
rect 395227 62485 397632 67323
rect 393531 62461 397632 62485
rect 388630 62448 397632 62461
rect 397882 62448 402258 67349
rect 402508 62448 406884 67349
rect 407134 62448 411510 67349
rect 411760 62448 416136 67349
rect 416386 62448 420762 67349
rect 421012 67324 425388 67349
rect 421012 62471 421550 67324
rect 422153 62471 425388 67324
rect 421012 62448 425388 62471
rect 425638 67316 430327 67349
rect 425638 62479 428531 67316
rect 429041 62479 430327 67316
rect 425638 62448 430327 62479
rect 282449 62444 430327 62448
rect 10930 62443 430327 62444
rect 430568 67346 439266 67349
rect 430568 67324 435109 67346
rect 430568 62472 431483 67324
rect 432140 62472 435109 67324
rect 430568 62462 435109 62472
rect 435349 62462 439266 67346
rect 430568 62448 439266 62462
rect 439516 62448 443892 67349
rect 444142 62448 448518 67349
rect 448768 62448 453044 67349
rect 453294 62448 457770 67349
rect 458020 62448 462196 67349
rect 462446 67277 471248 67349
rect 462446 62510 465312 67277
rect 467131 62510 471248 67277
rect 462446 62448 471248 62510
rect 471498 62448 476174 67349
rect 476424 62448 480900 67349
rect 481150 67346 494578 67349
rect 481150 67310 490841 67346
rect 481150 62481 486318 67310
rect 486562 67294 490841 67310
rect 486562 62510 487006 67294
rect 488459 62510 490841 67294
rect 486562 62481 490841 62510
rect 481150 62471 490841 62481
rect 491077 62471 494578 67346
rect 481150 62448 494578 62471
rect 494828 67291 500401 67349
rect 494828 62507 498357 67291
rect 499810 62507 500401 67291
rect 494828 62448 500401 62507
rect 430568 62445 500401 62448
rect 500662 67349 571358 67353
rect 500662 62448 503780 67349
rect 504030 67340 571358 67349
rect 504030 67325 571006 67340
rect 504030 67324 558449 67325
rect 504030 67281 529618 67324
rect 504030 67262 509143 67281
rect 504030 62478 505496 67262
rect 506949 62497 509143 67262
rect 510596 62497 516863 67281
rect 518316 62497 529618 67281
rect 506949 62478 529618 62497
rect 504030 62466 529618 62478
rect 529869 67322 558449 67324
rect 529869 62471 537554 67322
rect 537879 67296 558449 67322
rect 537879 62471 539787 67296
rect 529869 62466 539787 62471
rect 504030 62457 539787 62466
rect 540637 62481 558449 67296
rect 558832 67301 571006 67325
rect 558832 62481 562936 67301
rect 540637 62472 562936 62481
rect 563908 66204 571006 67301
rect 571316 66204 571358 67340
rect 563908 66142 571358 66204
rect 563908 62472 566431 66142
rect 540637 62457 566431 62472
rect 504030 62448 566431 62457
rect 500662 62445 566431 62448
rect 430568 62443 566431 62445
rect 10930 62390 566431 62443
rect 58920 61688 60140 62390
rect 414838 61829 415704 61941
rect 42688 61108 80338 61688
rect 290382 61397 344299 61438
rect 83814 61116 84680 61171
rect 83814 60071 83875 61116
rect 43451 59461 83875 60071
rect 83814 58740 83875 59461
rect 84621 58740 84680 61116
rect 290382 59454 290503 61397
rect 291181 60809 344299 61397
rect 291181 59454 291291 60809
rect 414838 60678 414932 61829
rect 415612 60678 415704 61829
rect 414838 60575 415704 60678
rect 290382 59409 291291 59454
rect 83814 58670 84680 58740
rect 415095 57822 415495 60575
rect 415095 57384 427817 57822
rect 415095 54589 415495 57384
rect 429227 56295 430088 56297
rect 415939 55885 430088 56295
rect 415095 54151 427764 54589
rect 347494 53468 391206 53534
rect 347494 53463 389744 53468
rect 347494 53453 382998 53463
rect 347494 51577 347668 53453
rect 350 51220 7234 51540
rect 347473 50652 347668 51577
rect 351477 50652 382998 53453
rect 347473 50614 382998 50652
rect 383893 50614 389744 53463
rect 347473 50582 389744 50614
rect 390995 50582 391206 53468
rect 429227 53031 430088 55885
rect 573027 55200 574600 55520
rect 570970 54200 574282 54520
rect 415939 52621 430088 53031
rect 0 50220 6247 50540
rect 347473 50534 391206 50582
rect 350 30220 7116 30540
rect 0 29220 6738 29540
rect -6 13157 8828 16557
rect 347473 15393 350473 50534
rect 429227 48534 430088 52621
rect 295413 15312 350473 15393
rect 295413 14892 339670 15312
rect 340952 14892 350473 15312
rect 295413 14786 350473 14892
rect 352971 48473 525803 48534
rect 352971 48413 405504 48473
rect 352971 45614 391494 48413
rect 392733 45614 405504 48413
rect 352971 45583 405504 45614
rect 406457 48410 525803 48473
rect 406457 45689 521477 48410
rect 525395 45689 525803 48410
rect 406457 45583 525803 45689
rect 352971 45534 525803 45583
rect 352971 23750 355971 45534
rect 368182 45515 369817 45534
rect 368182 44750 368294 45515
rect 369665 44750 369817 45515
rect 368182 44591 369817 44750
rect 374840 39680 385786 39726
rect 374840 39126 384400 39680
rect 385734 39126 385786 39680
rect 374840 39078 385786 39126
rect 373034 23750 373620 38182
rect 352971 22888 373620 23750
rect 374840 22898 375288 39078
rect -6 13072 82570 13157
rect -6 11629 81321 13072
rect 82276 11629 82570 13072
rect -6 11557 82570 11629
rect 295413 11968 296176 14786
rect 352971 13855 355971 22888
rect 373034 22104 373620 22888
rect 376786 22104 377372 38182
rect 378654 22898 379102 39078
rect 380598 22104 381184 38196
rect 382312 22946 382760 39078
rect 572442 34200 574600 34520
rect 571033 33200 574302 33520
rect 567335 27368 574604 30557
rect 469927 24357 488773 25957
rect 373034 21694 373732 22104
rect 376786 21694 377498 22104
rect 380598 21862 381264 22104
rect 380598 21694 381262 21862
rect 296867 13008 355971 13855
rect 358278 21284 371511 21597
rect 358278 20548 363198 21284
rect 363516 20548 371511 21284
rect 373034 21046 381262 21694
rect 358278 20414 371511 20548
rect 469927 20414 471527 24357
rect 358278 19997 471527 20414
rect 295413 11885 341089 11968
rect 295413 11465 339692 11885
rect 340974 11465 341089 11885
rect 295413 11361 341089 11465
rect 358278 9691 359878 19997
rect 132644 9650 359878 9691
rect -6 9553 8828 9557
rect -6 9464 84002 9553
rect -6 8021 82751 9464
rect 83706 8021 84002 9464
rect 132644 8142 132718 9650
rect 133480 8142 359878 9650
rect 132644 8091 359878 8142
rect 360678 18014 369111 19197
rect 369911 18814 471527 19997
rect 472435 21849 485794 23449
rect 472435 18014 474035 21849
rect 479014 20475 480562 20654
rect 475441 19695 476857 19700
rect 475434 19501 478564 19695
rect 475434 18455 475586 19501
rect 478387 18455 478564 19501
rect 475434 18311 478564 18455
rect 479014 18553 479182 20475
rect 480378 18553 480562 20475
rect 360678 17597 474035 18014
rect -6 7953 84002 8021
rect -6 4557 8828 7953
rect 360678 7291 362278 17597
rect 364507 16947 365371 17028
rect 364507 15024 364589 16947
rect 365295 15024 365371 16947
rect 363618 14724 364152 14764
rect 363618 13435 363655 14724
rect 364110 13435 364152 14724
rect 363618 10400 364152 13435
rect 364507 13158 365371 15024
rect 364507 11594 364566 13158
rect 365310 11594 365371 13158
rect 364507 11533 365371 11594
rect 365805 16970 366642 17055
rect 365805 15047 365875 16970
rect 366581 15047 366642 16970
rect 367511 16414 474035 17597
rect 363646 8230 364152 10400
rect 365805 11319 366642 15047
rect 365805 9755 365865 11319
rect 366609 9755 366642 11319
rect 365805 9697 366642 9755
rect 131408 7246 362278 7291
rect 131408 5738 131510 7246
rect 132272 5738 362278 7246
rect 131408 5691 362278 5738
rect 363618 4706 364152 8230
rect 475441 7697 476857 18311
rect 475441 6385 475597 7697
rect 476706 6385 476857 7697
rect 475441 6247 476857 6385
rect 479014 4706 480562 18553
rect 484194 8084 485794 21849
rect 487173 10906 488773 24357
rect 563945 25768 574604 27368
rect 563945 10906 565545 25768
rect 567335 25557 574604 25768
rect 567335 23553 574604 23557
rect 487173 10794 565545 10906
rect 487173 10414 487572 10794
rect 488240 10414 565545 10794
rect 487173 9306 565545 10414
rect 566768 18557 574604 23553
rect 566768 8084 568368 18557
rect 571842 16120 572162 16135
rect 571842 13520 572162 15800
rect 571842 13200 574600 13520
rect 572674 12200 574294 12520
rect 484194 6484 568368 8084
rect 90261 4673 514620 4706
rect 90261 4669 341501 4673
rect 90261 4664 338746 4669
rect 90261 4662 231731 4664
rect 90261 4661 173431 4662
rect 90261 4643 123625 4661
rect 90261 3174 91118 4643
rect 91406 3181 123625 4643
rect 123912 4622 173431 4661
rect 123912 3258 156181 4622
rect 157163 3258 173431 4622
rect 123912 3181 173431 3258
rect 91406 3176 173431 3181
rect 174106 4611 231731 4662
rect 174106 3227 215109 4611
rect 216072 3227 231731 4611
rect 174106 3176 231731 3227
rect 232396 4660 338746 4664
rect 232396 3198 254124 4660
rect 254704 4628 338746 4660
rect 254704 3262 277360 4628
rect 278170 4600 338746 4628
rect 278170 3262 286652 4600
rect 254704 3247 286652 3262
rect 287645 3247 338746 4600
rect 254704 3198 338746 3247
rect 232396 3176 338746 3198
rect 91406 3174 338746 3176
rect 90261 3172 338746 3174
rect 339105 3176 341501 4669
rect 341760 4638 514620 4673
rect 341760 4624 494902 4638
rect 341760 3276 490718 4624
rect 491898 3276 494902 4624
rect 341760 3202 494902 3276
rect 496002 4634 514620 4638
rect 496002 4588 513408 4634
rect 496002 3217 509316 4588
rect 510361 3217 513408 4588
rect 496002 3202 513408 3217
rect 341760 3198 513408 3202
rect 514508 3198 514620 4634
rect 341760 3176 514620 3198
rect 339105 3172 514620 3176
rect 90261 3138 514620 3172
rect 90261 2250 520026 2281
rect 90261 2245 230517 2250
rect 90261 2237 172217 2245
rect 90261 2234 124153 2237
rect 90261 765 90590 2234
rect 90878 765 124153 2234
rect 90261 757 124153 765
rect 124440 2183 172217 2237
rect 124440 819 148608 2183
rect 149590 819 172217 2183
rect 124440 759 172217 819
rect 172892 2191 230517 2245
rect 172892 807 207569 2191
rect 208532 807 230517 2191
rect 172892 759 230517 807
rect 231189 2237 520026 2250
rect 231189 2235 341930 2237
rect 231189 759 251034 2235
rect 124440 757 251034 759
rect 90261 751 251034 757
rect 251979 2213 341930 2235
rect 251979 786 279768 2213
rect 280605 2206 341930 2213
rect 280605 2173 294538 2206
rect 280605 820 288423 2173
rect 289416 820 294538 2173
rect 280605 796 294538 820
rect 294988 796 341930 2206
rect 280605 786 341930 796
rect 251979 751 341930 786
rect 90261 747 341930 751
rect 342210 2226 520026 2237
rect 342210 770 364588 2226
rect 365003 2210 520026 2226
rect 365003 2202 500288 2210
rect 365003 2136 485221 2202
rect 365003 824 475597 2136
rect 476706 843 485221 2136
rect 486580 843 500288 2202
rect 476706 824 500288 843
rect 365003 774 500288 824
rect 501388 2172 518780 2210
rect 501388 801 503942 2172
rect 504987 801 518780 2172
rect 501388 774 518780 801
rect 519880 774 520026 2210
rect 365003 770 520026 774
rect 342210 747 520026 770
rect 90261 713 520026 747
use analog_textblock  analog_textblock_0
timestamp 1731170561
transform 1 0 -308709 0 1 -83309
box 542248 94794 556139 108878
use cv3_via2_3cut  cv3_via2_3cut_0
timestamp 1719174692
transform 1 0 5246 0 1 1065
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_1
timestamp 1719174692
transform 1 0 4310 0 1 2600
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_2
timestamp 1719174692
transform 1 0 3826 0 1 2088
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_3
timestamp 1719174692
transform 1 0 4771 0 1 1574
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_4
timestamp 1719174692
transform 0 1 -50971 -1 0 542921
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_5
timestamp 1719174692
transform 0 1 -51081 -1 0 543267
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_6
timestamp 1719174692
transform 0 1 182599 -1 0 542922
box 542198 73062 542469 73190
use cv3_via2_3cut  cv3_via2_3cut_7
timestamp 1719174692
transform 0 1 182972 -1 0 543248
box 542198 73062 542469 73190
use cv3_via2_6cut  cv3_via2_6cut_0
timestamp 1719259570
transform 1 0 148608 0 1 75223
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_1
timestamp 1719259570
transform 1 0 144626 0 1 74711
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_2
timestamp 1719259570
transform 1 0 199710 0 1 70103
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_3
timestamp 1719259570
transform 1 0 204700 0 1 71639
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_4
timestamp 1719259570
transform 1 0 381802 0 1 75223
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_5
timestamp 1719259570
transform 1 0 375429 0 1 74711
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_6
timestamp 1719259570
transform 1 0 445726 0 1 73687
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_7
timestamp 1719259570
transform 1 0 436509 0 1 70103
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_8
timestamp 1719259570
transform 1 0 80667 0 1 64467
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_9
timestamp 1719259570
transform 1 0 127892 0 1 64983
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_10
timestamp 1719259570
transform 1 0 131589 0 1 69083
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_11
timestamp 1719259570
transform 1 0 225586 0 1 64476
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_12
timestamp 1719259570
transform 1 0 317159 0 1 67029
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_13
timestamp 1719259570
transform 1 0 316291 0 1 66515
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_14
timestamp 1719259570
transform 1 0 361425 0 1 67544
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_15
timestamp 1719259570
transform 1 0 360883 0 1 68057
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_16
timestamp 1719259570
transform 1 0 418789 0 1 61359
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_17
timestamp 1719259570
transform 1 0 404256 0 1 69084
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_18
timestamp 1719259570
transform 1 0 408781 0 1 68564
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_19
timestamp 1719259570
transform 1 0 402350 0 1 61365
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_20
timestamp 1719259570
transform 1 0 188172 0 1 63961
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_21
timestamp 1719259570
transform 1 0 468846 0 1 64984
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_22
timestamp 1719259570
transform 1 0 450364 0 1 64466
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_23
timestamp 1719259570
transform 1 0 190155 0 1 68558
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_24
timestamp 1719259570
transform 1 0 227636 0 1 64992
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_25
timestamp 1719259570
transform 1 0 211782 0 1 65486
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_26
timestamp 1719259570
transform 1 0 220834 0 1 70624
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_27
timestamp 1719259570
transform 1 0 216322 0 1 71632
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_28
timestamp 1719259570
transform 1 0 236774 0 1 71128
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_29
timestamp 1719259570
transform 1 0 241262 0 1 66002
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_30
timestamp 1719259570
transform 1 0 232264 0 1 72164
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_31
timestamp 1719259570
transform 1 0 454918 0 1 73704
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_32
timestamp 1719259570
transform 1 0 464312 0 1 67548
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_33
timestamp 1719259570
transform 1 0 482726 0 1 73178
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_34
timestamp 1719259570
transform 1 0 491984 0 1 67034
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_35
timestamp 1719259570
transform 1 0 487371 0 1 68065
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_36
timestamp 1719259570
transform 1 0 166897 0 1 62939
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_37
timestamp 1719259570
transform 1 0 225857 0 1 63451
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_38
timestamp 1719259570
transform 1 0 286788 0 1 68568
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_39
timestamp 1719259570
transform 1 0 286948 0 1 61908
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_40
timestamp 1719259570
transform 1 0 287144 0 1 69081
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_41
timestamp 1719259570
transform 1 0 287447 0 1 62422
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_42
timestamp 1719259570
transform 1 0 189501 0 1 66008
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_43
timestamp 1719259570
transform 1 0 130802 0 1 65497
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_44
timestamp 1719259570
transform 1 0 143964 0 1 70615
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_45
timestamp 1719259570
transform 1 0 204239 0 1 69591
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_46
timestamp 1719259570
transform 1 0 371915 0 1 72663
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_47
timestamp 1719259570
transform 1 0 441203 0 1 69591
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_50
timestamp 1719259570
transform 1 0 468890 0 1 66530
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_62
timestamp 1719259570
transform 1 0 459618 0 1 72656
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_68
timestamp 1719259570
transform 1 0 473518 0 1 64982
box 3030 432 3561 574
use cv3_via2_6cut  cv3_via2_6cut_73
timestamp 1719259570
transform 1 0 478144 0 1 74200
box 3030 432 3561 574
use cv3_via2_8cut  cv3_via2_8cut_0
timestamp 1719106786
transform 0 1 -13629 -1 0 68640
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_1
timestamp 1719106786
transform 0 1 -9635 -1 0 69033
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_2
timestamp 1719106786
transform 1 0 565604 0 1 4054
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_3
timestamp 1719106786
transform 1 0 -1180 0 1 3618
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_4
timestamp 1719106786
transform 1 0 -1780 0 1 4146
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_5
timestamp 1719106786
transform 1 0 -2368 0 1 4646
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_6
timestamp 1719106786
transform 1 0 -2962 0 1 5174
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_7
timestamp 1719106786
transform 1 0 -3550 0 1 5662
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_8
timestamp 1719106786
transform 1 0 -4142 0 1 6180
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_9
timestamp 1719106786
transform 1 0 563076 0 1 4060
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_10
timestamp 1719106786
transform 1 0 563716 0 1 4058
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_11
timestamp 1719106786
transform 1 0 564342 0 1 4058
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_12
timestamp 1719106786
transform 1 0 564976 0 1 4058
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_13
timestamp 1719106786
transform 1 0 81643 0 1 30693
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_14
timestamp 1719106786
transform 1 0 186486 0 1 -14153
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_15
timestamp 1719106786
transform 1 0 127148 0 1 -27662
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_16
timestamp 1719106786
transform 0 1 112197 -1 0 40498
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_17
timestamp 1719106786
transform 0 1 169327 -1 0 40649
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_18
timestamp 1719106786
transform 1 0 185837 0 1 -27526
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_30
timestamp 1719106786
transform 0 1 -35190 -1 0 108430
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_31
timestamp 1719106786
transform 0 1 -44832 -1 0 109328
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_32
timestamp 1719106786
transform 0 1 -40010 -1 0 108724
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_33
timestamp 1719106786
transform 0 1 -20668 -1 0 102553
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_34
timestamp 1719106786
transform 0 1 -30352 -1 0 103486
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_35
timestamp 1719106786
transform 0 1 -25472 -1 0 102843
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_36
timestamp 1719106786
transform 1 0 -1186 0 1 39024
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_37
timestamp 1719106786
transform 1 0 -1782 0 1 33170
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_38
timestamp 1719106786
transform 1 0 -2366 0 1 39330
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_39
timestamp 1719106786
transform 1 0 -3554 0 1 40120
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_40
timestamp 1719106786
transform 1 0 -4142 0 1 34276
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_41
timestamp 1719106786
transform 1 0 -2962 0 1 33468
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_43
timestamp 1719106786
transform 0 1 112197 -1 0 40138
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_45
timestamp 1719106786
transform 1 0 248810 0 1 -38531
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_47
timestamp 1719106786
transform 0 1 169327 -1 0 40289
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_48
timestamp 1719106786
transform 1 0 249184 0 1 -38716
box 6850 62208 6998 62544
use cv3_via2_9cut  cv3_via2_9cut_0
timestamp 1719106980
transform 1 0 3778 0 1 -4572
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_2
timestamp 1719106980
transform 1 0 1884 0 1 -3040
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_6
timestamp 1719106980
transform 1 0 3154 0 1 -4056
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_7
timestamp 1719106980
transform 1 0 -219670 0 1 -470
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_8
timestamp 1719106980
transform 1 0 -225294 0 1 -4576
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_9
timestamp 1719106980
transform 1 0 -224798 0 1 -4060
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_10
timestamp 1719106980
transform 1 0 -224274 0 1 -3544
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_11
timestamp 1719106980
transform 1 0 -223758 0 1 -3028
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_12
timestamp 1719106980
transform 1 0 -223248 0 1 -2518
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_13
timestamp 1719106980
transform 1 0 -222732 0 1 -1492
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_14
timestamp 1719106980
transform 1 0 -222236 0 1 -2016
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_15
timestamp 1719106980
transform 1 0 -221706 0 1 2604
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_16
timestamp 1719106980
transform 1 0 -221210 0 1 2088
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_17
timestamp 1719106980
transform 1 0 -217106 0 1 1572
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_18
timestamp 1719106980
transform 1 0 -217628 0 1 1064
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_19
timestamp 1719106980
transform 1 0 -218120 0 1 544
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_20
timestamp 1719106980
transform 1 0 -218642 0 1 36
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_21
timestamp 1719106980
transform 1 0 -219154 0 1 -980
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_36
timestamp 1719106980
transform 1 0 -286370 0 1 8746
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_37
timestamp 1719106980
transform 1 0 -331132 0 1 -1504
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_38
timestamp 1719106980
transform 1 0 -290490 0 1 8230
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_39
timestamp 1719106980
transform 1 0 -290890 0 1 6696
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_40
timestamp 1719106980
transform 1 0 -295016 0 1 6184
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_41
timestamp 1719106980
transform 1 0 -295410 0 1 7720
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_42
timestamp 1719106980
transform 1 0 -299526 0 1 7204
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_43
timestamp 1719106980
transform 1 0 -299932 0 1 4646
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_44
timestamp 1719106980
transform 1 0 -304056 0 1 4138
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_45
timestamp 1719106980
transform 1 0 -304450 0 1 5676
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_46
timestamp 1719106980
transform 1 0 -308564 0 1 5162
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_47
timestamp 1719106980
transform 1 0 -308960 0 1 3622
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_48
timestamp 1719106980
transform 1 0 -313072 0 1 3114
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_49
timestamp 1719106980
transform 1 0 -313472 0 1 1063
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_50
timestamp 1719106980
transform 1 0 -317596 0 1 1569
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_51
timestamp 1719106980
transform 1 0 -317996 0 1 37
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_52
timestamp 1719106980
transform 1 0 -322104 0 1 548
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_53
timestamp 1719106980
transform 1 0 -322506 0 1 -982
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_54
timestamp 1719106980
transform 1 0 -326620 0 1 -470
box 568286 66860 568540 67110
use cv3_via2_9cut  cv3_via2_9cut_55
timestamp 1719106980
transform 1 0 -327018 0 1 -2004
box 568286 66860 568540 67110
use cv3_via2_36cut  cv3_via2_36cut_0
timestamp 1719173892
transform 1 0 3800 0 1 2600
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_1
timestamp 1719173892
transform 1 0 11843 0 1 2078
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_2
timestamp 1719173892
transform -1 0 1101612 0 -1 173009
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_3
timestamp 1719173892
transform 1 0 11844 0 1 -11762
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_4
timestamp 1719173892
transform 1 0 -4370 0 1 -31390
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_5
timestamp 1719173892
transform 1 0 3992 0 1 -32459
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_6
timestamp 1719173892
transform 1 0 -4050 0 1 -43797
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_7
timestamp 1719173892
transform 1 0 3994 0 1 -40590
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_8
timestamp 1719173892
transform 1 0 -4900 0 1 -45623
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_9
timestamp 1719173892
transform 1 0 3143 0 1 -47939
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_10
timestamp 1719173892
transform 1 0 -4900 0 1 -57058
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_11
timestamp 1719173892
transform 1 0 3144 0 1 -58186
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_12
timestamp 1719173892
transform 1 0 -5200 0 1 -58970
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_13
timestamp 1719173892
transform 1 0 2872 0 1 -64495
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_14
timestamp 1719173892
transform 1 0 -611 0 1 -58515
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_15
timestamp 1719173892
transform 1 0 2844 0 1 -72102
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_16
timestamp 1719173892
transform 1 0 -8654 0 1 -72094
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_17
timestamp 1719173892
transform 1 0 -616 0 1 -72082
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_18
timestamp 1719173892
transform 1 0 -5200 0 1 -71489
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_19
timestamp 1719173892
transform 0 1 -47585 -1 0 652338
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_20
timestamp 1719173892
transform 0 1 -48085 -1 0 658204
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_21
timestamp 1719173892
transform 0 1 -48688 -1 0 664064
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_22
timestamp 1719173892
transform 1 0 -20498 0 1 -71679
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_23
timestamp 1719173892
transform 1 0 -8659 0 1 -59061
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_24
timestamp 1719173892
transform 1 0 -8365 0 1 -58058
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_25
timestamp 1719173892
transform 1 0 -333 0 1 -58107
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_26
timestamp 1719173892
transform 1 0 -7501 0 1 -32421
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_27
timestamp 1719173892
transform 1 0 -8365 0 1 -45615
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_28
timestamp 1719173892
transform 1 0 -7506 0 1 -44736
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_29
timestamp 1719173892
transform 1 0 -452048 0 1 22210
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_30
timestamp 1719173892
transform 1 0 -317 0 1 -45183
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_31
timestamp 1719173892
transform 1 0 539 0 1 -44800
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_32
timestamp 1719173892
transform 1 0 523 0 1 -32169
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_33
timestamp 1719173892
transform 1 0 -453854 0 1 21800
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_34
timestamp 1719173892
transform 1 0 -464270 0 1 21415
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_35
timestamp 1719173892
transform 1 0 -467066 0 1 18882
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_36
timestamp 1719173892
transform 1 0 -63730 0 1 19490
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_37
timestamp 1719173892
transform 1 0 -47954 0 1 20110
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_38
timestamp 1719173892
transform 1 0 -49682 0 1 21759
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_39
timestamp 1719173892
transform 1 0 -62568 0 1 21506
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_40
timestamp 1719173892
transform 1 0 -465468 0 1 19482
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_41
timestamp 1719173892
transform 1 0 -466582 0 1 21008
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_42
timestamp 1719173892
transform 1 0 -450886 0 1 17014
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_43
timestamp 1719173892
transform 1 0 -452674 0 1 17602
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_44
timestamp 1719173892
transform 1 0 -277174 0 1 21530
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_45
timestamp 1719173892
transform 1 0 -290766 0 1 19498
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_46
timestamp 1719173892
transform 1 0 -291550 0 1 20756
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_47
timestamp 1719173892
transform 1 0 -327175 0 1 14880
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_48
timestamp 1719173892
transform 1 0 -290230 0 1 21126
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_49
timestamp 1719173892
transform 1 0 -275592 0 1 21932
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_50
timestamp 1719173892
transform 1 0 -274390 0 1 18266
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_51
timestamp 1719173892
transform 1 0 -276074 0 1 17648
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_52
timestamp 1719173892
transform 1 0 -242340 0 1 19510
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_53
timestamp 1719173892
transform 1 0 -244194 0 1 18878
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_54
timestamp 1719173892
transform 0 1 171756 -1 0 654774
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_55
timestamp 1719173892
transform 1 0 -227398 0 1 17652
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_56
timestamp 1719173892
transform 1 0 -64096 0 1 22056
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_57
timestamp 1719173892
transform 1 0 -91900 0 1 15187
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_58
timestamp 1719173892
transform 1 0 -49632 0 1 17612
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_59
timestamp 1719173892
transform 1 0 -48518 0 1 21294
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_60
timestamp 1719173892
transform 1 0 -527874 0 1 -72782
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_61
timestamp 1719173892
transform 1 0 -539378 0 1 -73970
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_62
timestamp 1719173892
transform 1 0 -535932 0 1 -72190
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_63
timestamp 1719173892
transform 1 0 -531344 0 1 -73384
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_64
timestamp 1719173892
transform 1 0 -539386 0 1 -59376
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_65
timestamp 1719173892
transform 1 0 -539382 0 1 -56546
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_66
timestamp 1719173892
transform 1 0 -535938 0 1 -58934
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_67
timestamp 1719173892
transform 1 0 -531354 0 1 -57622
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_68
timestamp 1719173892
transform 1 0 -535938 0 1 -44934
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_69
timestamp 1719173892
transform 1 0 -539394 0 1 -42538
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_70
timestamp 1719173892
transform 1 0 -539372 0 1 -45374
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_71
timestamp 1719173892
transform 1 0 -531338 0 1 -43638
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_72
timestamp 1719173892
transform 1 0 -539378 0 1 -31478
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_73
timestamp 1719173892
transform 1 0 -527892 0 1 -30632
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_74
timestamp 1719173892
transform 1 0 -536082 0 1 -15524
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_75
timestamp 1719173892
transform 1 0 -539540 0 1 -14322
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_76
timestamp 1719173892
transform 1 0 -531498 0 1 -2854
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_77
timestamp 1719173892
transform 1 0 -528048 0 1 -2208
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_78
timestamp 1719173892
transform 1 0 -527892 0 1 -58632
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_79
timestamp 1719173892
transform 1 0 -531348 0 1 -58990
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_80
timestamp 1719173892
transform -1 0 569655 0 -1 188591
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_81
timestamp 1719173892
transform -1 0 570526 0 -1 200359
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_82
timestamp 1719173892
transform 1 0 -527876 0 1 -58042
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_83
timestamp 1719173892
transform -1 0 570167 0 -1 194464
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_84
timestamp 1719173892
transform 1 0 -535936 0 1 -57616
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_85
timestamp 1719173892
transform 1 0 -62448 0 1 -84652
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_86
timestamp 1719173892
transform 1 0 -243278 0 1 22246
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_87
timestamp 1719173892
transform 1 0 -527892 0 1 -44632
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_88
timestamp 1719173892
transform 1 0 -531340 0 1 -45030
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_89
timestamp 1719173892
transform 1 0 -241112 0 1 21772
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_90
timestamp 1719173892
transform 1 0 -527876 0 1 -44042
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_91
timestamp 1719173892
transform 1 0 -227852 0 1 21394
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_92
timestamp 1719173892
transform 1 0 -535936 0 1 -43616
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_93
timestamp 1719173892
transform 1 0 -226182 0 1 20952
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_94
timestamp 1719173892
transform 1 0 -535938 0 1 -30934
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_95
timestamp 1719173892
transform 1 0 -531342 0 1 -31092
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_96
timestamp 1719173892
transform 0 1 414496 -1 0 654500
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_97
timestamp 1719173892
transform 0 1 445030 -1 0 635633
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_98
timestamp 1719173892
transform 1 0 -528044 0 1 -15942
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_99
timestamp 1719173892
transform 1 0 -531506 0 1 -15474
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_100
timestamp 1719173892
transform 1 0 -536088 0 1 -2764
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_101
timestamp 1719173892
transform 1 0 -539542 0 1 -3242
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_102
timestamp 1719173892
transform 0 1 434517 -1 0 636083
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_103
timestamp 1719173892
transform -1 0 609378 0 -1 170102
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_104
timestamp 1719173892
transform 0 1 479223 -1 0 564587
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_105
timestamp 1719173892
transform 0 1 -1208 -1 0 661816
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_106
timestamp 1719173892
transform 0 1 251270 -1 0 612686
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_107
timestamp 1719173892
transform 0 1 258956 -1 0 615184
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_108
timestamp 1719173892
transform 0 1 258444 -1 0 614888
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_109
timestamp 1719173892
transform 0 1 257922 -1 0 614582
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_110
timestamp 1719173892
transform 0 1 257414 -1 0 614290
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_111
timestamp 1719173892
transform 0 1 256912 -1 0 613988
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_112
timestamp 1719173892
transform 0 1 256386 -1 0 613690
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_113
timestamp 1719173892
transform 0 1 -17906 -1 0 632403
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_114
timestamp 1719173892
transform 1 0 -541654 0 1 20114
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_115
timestamp 1719173892
transform 0 1 254858 -1 0 614796
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_116
timestamp 1719173892
transform 0 1 254350 -1 0 614498
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_117
timestamp 1719173892
transform 0 1 253828 -1 0 614188
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_118
timestamp 1719173892
transform 0 1 253308 -1 0 613890
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_119
timestamp 1719173892
transform 0 1 252802 -1 0 613594
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_120
timestamp 1719173892
transform 0 1 252284 -1 0 613296
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_121
timestamp 1719173892
transform 0 1 251772 -1 0 612992
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_122
timestamp 1719173892
transform 0 1 250752 -1 0 612400
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_123
timestamp 1719173892
transform 1 0 -542066 0 1 19490
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_124
timestamp 1719173892
transform 1 0 -512452 0 1 17018
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_125
timestamp 1719173892
transform 1 0 -511322 0 1 18870
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_126
timestamp 1719173892
transform 1 0 -511840 0 1 17646
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_127
timestamp 1719173892
transform 1 0 -542554 0 1 18254
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_128
timestamp 1719173892
transform 0 1 -27645 -1 0 632520
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_129
timestamp 1719173892
transform 0 1 -7121 -1 0 632357
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_130
timestamp 1719173892
transform 1 0 8402 0 1 -10627
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_131
timestamp 1719173892
transform 1 0 3800 0 1 -11007
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_132
timestamp 1719173892
transform 1 0 359 0 1 -10710
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_133
timestamp 1719173892
transform 1 0 -261490 0 1 20134
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_134
timestamp 1719173892
transform 1 0 -262734 0 1 18878
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_135
timestamp 1719173892
transform 1 0 -255560 0 1 19518
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_136
timestamp 1719173892
transform 1 0 -249646 0 1 18258
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_137
timestamp 1719173892
transform 1 0 -256788 0 1 17628
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_138
timestamp 1719173892
transform 1 0 -250908 0 1 16996
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_139
timestamp 1719173892
transform 0 1 453807 -1 0 634700
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_140
timestamp 1719173892
transform -1 0 1107089 0 -1 188198
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_141
timestamp 1719173892
transform 1 0 -278402 0 1 -72872
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_142
timestamp 1719173892
transform 1 0 -274932 0 1 -72872
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_143
timestamp 1719173892
transform 1 0 -274974 0 1 -59780
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_144
timestamp 1719173892
transform 1 0 -278402 0 1 -59832
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_145
timestamp 1719173892
transform 0 1 455292 -1 0 633687
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_146
timestamp 1719173892
transform 0 1 454746 -1 0 634072
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_147
timestamp 1719173892
transform 1 0 -225482 0 1 18252
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_148
timestamp 1719173892
transform 0 1 236872 -1 0 654564
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_149
timestamp 1719173892
transform 0 1 235168 -1 0 662598
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_150
timestamp 1719173892
transform 0 1 221980 -1 0 662620
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_151
timestamp 1719173892
transform 0 1 220152 -1 0 654564
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_152
timestamp 1719173892
transform 0 1 188056 -1 0 654668
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_153
timestamp 1719173892
transform 0 1 186520 -1 0 662746
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_154
timestamp 1719173892
transform 0 1 173396 -1 0 662766
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_155
timestamp 1719173892
transform 0 1 400416 -1 0 662576
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_156
timestamp 1719173892
transform 0 1 398922 -1 0 654522
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_157
timestamp 1719173892
transform 0 1 -2736 -1 0 654106
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_158
timestamp 1719173892
transform 0 1 413604 -1 0 662556
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_159
timestamp 1719173892
transform 0 1 415566 -1 0 640527
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_160
timestamp 1719173892
transform 0 1 11648 -1 0 654084
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_161
timestamp 1719173892
transform 0 1 10644 -1 0 662232
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_162
timestamp 1719173892
transform 0 1 -544 -1 0 663560
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_163
timestamp 1719173892
transform 1 0 262 0 1 -30958
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_164
timestamp 1719173892
transform 0 1 479869 -1 0 564196
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_165
timestamp 1719173892
transform 0 1 478040 -1 0 565728
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_166
timestamp 1719173892
transform 1 0 9532 0 1 -30502
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_167
timestamp 1719173892
transform 0 1 437860 -1 0 611006
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_168
timestamp 1719173892
transform 0 1 449422 -1 0 610992
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_169
timestamp 1719173892
transform 0 1 449365 -1 0 607527
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_170
timestamp 1719173892
transform 0 1 437894 -1 0 607546
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_171
timestamp 1719173892
transform 0 1 454292 -1 0 634447
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_172
timestamp 1719173892
transform 1 0 -17021 0 1 -58286
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_173
timestamp 1719173892
transform 1 0 -17019 0 1 -45080
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_174
timestamp 1719173892
transform 1 0 -20482 0 1 -44540
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_175
timestamp 1719173892
transform 1 0 -20501 0 1 -58972
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_176
timestamp 1719173892
transform 1 0 -20471 0 1 -57886
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_177
timestamp 1719173892
transform 1 0 -16864 0 1 -75509
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_178
timestamp 1719173892
transform 1 0 -467557 0 1 17009
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_179
timestamp 1719173892
transform 1 0 -4195 0 1 20514
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_180
timestamp 1719173892
transform 1 0 -65406 0 1 18870
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_181
timestamp 1719173892
transform 1 0 -91923 0 1 18867
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_182
timestamp 1719173892
transform 1 0 -429349 0 1 14617
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_183
timestamp 1719173892
transform 1 0 -429341 0 1 18250
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_184
timestamp 1719173892
transform 1 0 -292690 0 1 18884
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_185
timestamp 1719173892
transform 1 0 -327194 0 1 17625
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_186
timestamp 1719173892
transform 1 0 -195027 0 1 15146
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_187
timestamp 1719173892
transform 1 0 -194976 0 1 19502
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_188
timestamp 1719173892
transform 0 1 86017 -1 0 635894
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_189
timestamp 1719173892
transform 1 0 -379587 0 1 18261
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_190
timestamp 1719173892
transform 1 0 -377121 0 1 17625
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_191
timestamp 1719173892
transform 0 1 64604 -1 0 636025
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_192
timestamp 1719173892
transform 0 1 83744 -1 0 661993
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_193
timestamp 1719173892
transform 0 1 86213 -1 0 661932
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_194
timestamp 1719173892
transform 0 1 83901 -1 0 635860
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_195
timestamp 1719173892
transform 0 1 86004 -1 0 643673
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_196
timestamp 1719173892
transform 0 1 83905 -1 0 643675
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_197
timestamp 1719173892
transform -1 0 711553 0 -1 186203
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_198
timestamp 1719173892
transform 0 -1 290881 -1 0 636009
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_199
timestamp 1719173892
transform 0 -1 288963 -1 0 652188
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_200
timestamp 1719173892
transform 0 1 297226 -1 0 635616
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_201
timestamp 1719173892
transform 0 1 300315 -1 0 651753
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_202
timestamp 1719173892
transform 0 1 320217 -1 0 635494
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_203
timestamp 1719173892
transform 0 1 318101 -1 0 635460
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_204
timestamp 1719173892
transform 0 1 320211 -1 0 643160
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_205
timestamp 1719173892
transform 0 1 318105 -1 0 643225
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_206
timestamp 1719173892
transform 0 1 320413 -1 0 661532
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_207
timestamp 1719173892
transform 0 1 317944 -1 0 661593
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_208
timestamp 1719173892
transform 0 -1 527809 -1 0 635627
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_209
timestamp 1719173892
transform 0 -1 523163 -1 0 651693
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_210
timestamp 1719173892
transform 1 0 -142925 0 1 18891
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_211
timestamp 1719173892
transform 1 0 -145409 0 1 19502
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_212
timestamp 1719173892
transform 0 1 65715 -1 0 652203
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_213
timestamp 1719173892
transform 1 0 -356541 0 -1 186463
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_214
timestamp 1719173892
transform -1 0 945923 0 -1 186693
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_215
timestamp 1719173892
transform 1 0 -121371 0 -1 186723
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_216
timestamp 1719173892
transform 0 1 459971 -1 0 640461
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_217
timestamp 1719173892
transform 0 1 459527 -1 0 640421
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_220
timestamp 1719173892
transform -1 0 876552 0 -1 152470
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_221
timestamp 1719173892
transform -1 0 874951 0 -1 152443
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_222
timestamp 1719173892
transform 1 0 -133419 0 1 -47639
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_223
timestamp 1719173892
transform 1 0 -162625 0 1 -48017
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_224
timestamp 1719173892
transform 1 0 -139036 0 1 -48028
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_225
timestamp 1719173892
transform 1 0 -119549 0 1 -47621
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_226
timestamp 1719173892
transform 1 0 -72362 0 1 -47981
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_227
timestamp 1719173892
transform 1 0 -71698 0 1 -30534
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_230
timestamp 1719173892
transform 1 0 -163363 0 1 -31660
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_231
timestamp 1719173892
transform 1 0 -369282 0 1 -30704
box 555256 92202 556228 92502
use cv3_via3_10cut  cv3_via3_10cut_0
timestamp 1719433677
transform 1 0 739 0 1 4137
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_1
timestamp 1719433677
transform 1 0 -349 0 1 3630
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_2
timestamp 1719433677
transform 1 0 -41458 0 1 3102
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_3
timestamp 1719433677
transform 1 0 -39867 0 1 2600
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_4
timestamp 1719433677
transform 1 0 -234437 0 1 2088
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_5
timestamp 1719433677
transform 1 0 -235482 0 1 1579
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_6
timestamp 1719433677
transform 1 0 -275438 0 1 1064
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_7
timestamp 1719433677
transform 1 0 -274321 0 1 553
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_8
timestamp 1719433677
transform 1 0 -357630 0 1 36
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_9
timestamp 1719433677
transform 1 0 -346738 0 1 -474
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_10
timestamp 1719433677
transform 1 0 105395 0 1 5169
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_11
timestamp 1719433677
transform 1 0 43869 0 1 -15339
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_12
timestamp 1719433677
transform 1 0 -399604 0 1 2598
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_13
timestamp 1719433677
transform 1 0 -399184 0 1 3112
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_14
timestamp 1719433677
transform 1 0 -399996 0 1 2088
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_15
timestamp 1719433677
transform 1 0 -400398 0 1 1578
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_16
timestamp 1719433677
transform 1 0 -398366 0 1 38
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_17
timestamp 1719433677
transform 1 0 -398860 0 1 -476
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_18
timestamp 1719433677
transform 1 0 -399264 0 1 -1996
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_19
timestamp 1719433677
transform 1 0 -399642 0 1 -2526
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_20
timestamp 1719433677
transform 1 0 -400054 0 1 -3040
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_21
timestamp 1719433677
transform 1 0 -400474 0 1 -3538
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_22
timestamp 1719433677
transform 1 0 -400850 0 1 -4054
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_23
timestamp 1719433677
transform 1 0 -401197 0 1 -4566
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_24
timestamp 1719433677
transform 1 0 -397966 0 1 554
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_25
timestamp 1719433677
transform 1 0 -396860 0 1 1066
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_26
timestamp 1719433677
transform 1 0 110389 0 1 -37340
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_27
timestamp 1719433677
transform 0 -1 613437 1 0 -397679
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_28
timestamp 1719433677
transform 0 -1 612659 1 0 -398334
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_29
timestamp 1719433677
transform 0 -1 613180 1 0 -398029
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_30
timestamp 1719433677
transform 1 0 111397 0 1 -23794
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_31
timestamp 1719433677
transform 0 1 473323 -1 0 480471
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_32
timestamp 1719433677
transform 0 1 472556 -1 0 479933
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_33
timestamp 1719433677
transform 0 1 473074 -1 0 480211
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_34
timestamp 1719433677
transform 1 0 112418 0 1 -10672
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_35
timestamp 1719433677
transform 0 1 473580 -1 0 493044
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_36
timestamp 1719433677
transform 1 0 111141 0 1 -2014
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_37
timestamp 1719433677
transform 1 0 112422 0 1 -4565
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_38
timestamp 1719433677
transform 1 0 112167 0 1 -4056
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_39
timestamp 1719433677
transform 1 0 111920 0 1 -3539
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_40
timestamp 1719433677
transform 1 0 111654 0 1 -3030
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_41
timestamp 1719433677
transform 1 0 111407 0 1 -2520
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_42
timestamp 1719433677
transform 1 0 110119 0 1 3109
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_43
timestamp 1719433677
transform 1 0 110886 0 1 1573
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_44
timestamp 1719433677
transform 1 0 110624 0 1 2090
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_45
timestamp 1719433677
transform 1 0 110370 0 1 2606
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_46
timestamp 1719433677
transform 1 0 -424442 0 1 -1752
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_47
timestamp 1719433677
transform 1 0 -424442 0 1 -4824
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_48
timestamp 1719433677
transform 1 0 -424442 0 1 -4312
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_49
timestamp 1719433677
transform 1 0 -424442 0 1 -3800
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_50
timestamp 1719433677
transform 1 0 -424442 0 1 -3288
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_51
timestamp 1719433677
transform 1 0 -424442 0 1 -2776
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_52
timestamp 1719433677
transform 1 0 -424442 0 1 -2264
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_53
timestamp 1719433677
transform 0 1 285226 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_54
timestamp 1719433677
transform 0 1 284202 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_55
timestamp 1719433677
transform 0 1 284714 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_56
timestamp 1719433677
transform 0 1 292394 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_57
timestamp 1719433677
transform 0 1 285738 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_58
timestamp 1719433677
transform 0 1 286250 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_59
timestamp 1719433677
transform 0 1 286762 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_60
timestamp 1719433677
transform 0 1 287274 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_61
timestamp 1719433677
transform 0 1 287786 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_62
timestamp 1719433677
transform 0 1 288298 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_63
timestamp 1719433677
transform 0 1 288810 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_64
timestamp 1719433677
transform 0 1 289322 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_65
timestamp 1719433677
transform 0 1 289834 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_66
timestamp 1719433677
transform 0 1 290346 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_67
timestamp 1719433677
transform 0 1 290858 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_68
timestamp 1719433677
transform 0 1 291370 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_69
timestamp 1719433677
transform 0 1 291882 -1 0 491549
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_70
timestamp 1719433677
transform 1 0 -180922 0 1 -69352
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_71
timestamp 1719433677
transform 1 0 -180923 0 1 -62619
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_72
timestamp 1719433677
transform 1 0 -180925 0 1 -63241
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_73
timestamp 1719433677
transform 1 0 -180923 0 1 -65109
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_74
timestamp 1719433677
transform 1 0 -180922 0 1 -70255
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_75
timestamp 1719433677
transform 1 0 -180925 0 1 -63859
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_76
timestamp 1719433677
transform 1 0 -180921 0 1 -64485
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_77
timestamp 1719433677
transform 0 1 214810 -1 0 491493
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_78
timestamp 1719433677
transform 0 1 211774 -1 0 491493
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_79
timestamp 1719433677
transform 0 1 213186 -1 0 491493
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_80
timestamp 1719433677
transform 0 1 213998 -1 0 491493
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_81
timestamp 1719433677
transform 0 1 215622 -1 0 491493
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_82
timestamp 1719433677
transform 0 1 212374 -1 0 491493
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_83
timestamp 1719433677
transform 1 0 107801 0 1 -728
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_84
timestamp 1719433677
transform 1 0 107801 0 1 5416
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_85
timestamp 1719433677
transform 1 0 107801 0 1 4904
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_86
timestamp 1719433677
transform 1 0 107801 0 1 4392
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_87
timestamp 1719433677
transform 1 0 107801 0 1 3880
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_88
timestamp 1719433677
transform 1 0 107801 0 1 3368
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_89
timestamp 1719433677
transform 1 0 107801 0 1 2856
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_90
timestamp 1719433677
transform 1 0 107801 0 1 2344
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_91
timestamp 1719433677
transform 1 0 107801 0 1 1832
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_92
timestamp 1719433677
transform 1 0 107801 0 1 1320
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_93
timestamp 1719433677
transform 1 0 107801 0 1 808
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_94
timestamp 1719433677
transform 1 0 107801 0 1 296
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_95
timestamp 1719433677
transform 1 0 107801 0 1 -216
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_96
timestamp 1719433677
transform 1 0 107801 0 1 -8408
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_97
timestamp 1719433677
transform 1 0 107801 0 1 -6360
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_98
timestamp 1719433677
transform 1 0 107801 0 1 -6872
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_99
timestamp 1719433677
transform 1 0 107801 0 1 -7384
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_100
timestamp 1719433677
transform 1 0 107801 0 1 -7896
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_101
timestamp 1719433677
transform 1 0 -350550 0 1 -30556
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_102
timestamp 1719433677
transform 1 0 -350552 0 1 -24494
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_103
timestamp 1719433677
transform 1 0 12242 0 1 -1240
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_104
timestamp 1719433677
transform 1 0 12244 0 1 -5846
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_105
timestamp 1719433677
transform 1 0 12236 0 1 -5332
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_106
timestamp 1719433677
transform 1 0 -173599 0 1 38482
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_107
timestamp 1719433677
transform 1 0 -173599 0 1 42214
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_108
timestamp 1719433677
transform 1 0 -173599 0 1 41592
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_109
timestamp 1719433677
transform 1 0 -173599 0 1 40970
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_110
timestamp 1719433677
transform 1 0 -173599 0 1 40348
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_111
timestamp 1719433677
transform 1 0 -173599 0 1 39726
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_112
timestamp 1719433677
transform 1 0 -173599 0 1 39104
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_113
timestamp 1719433677
transform 1 0 94352 0 1 -6616
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_114
timestamp 1719433677
transform 0 1 283178 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_115
timestamp 1719433677
transform 1 0 -367686 0 1 -7124
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_116
timestamp 1719433677
transform 1 0 -367704 0 1 3904
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_117
timestamp 1719433677
transform 0 1 275498 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_118
timestamp 1719433677
transform 0 1 276010 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_119
timestamp 1719433677
transform 0 1 276522 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_120
timestamp 1719433677
transform 0 1 277034 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_121
timestamp 1719433677
transform 0 1 277546 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_122
timestamp 1719433677
transform 0 1 278058 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_123
timestamp 1719433677
transform 0 1 278570 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_124
timestamp 1719433677
transform 0 1 279082 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_125
timestamp 1719433677
transform 0 1 279594 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_126
timestamp 1719433677
transform 0 1 280106 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_127
timestamp 1719433677
transform 0 1 280618 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_128
timestamp 1719433677
transform 0 1 281130 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_129
timestamp 1719433677
transform 0 1 281642 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_130
timestamp 1719433677
transform 0 1 282154 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_131
timestamp 1719433677
transform 0 1 282666 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_132
timestamp 1719433677
transform 0 1 284202 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_133
timestamp 1719433677
transform 0 1 283690 -1 0 439816
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_134
timestamp 1719433677
transform 1 0 -257952 0 1 42216
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_135
timestamp 1719433677
transform 1 0 -209928 0 1 42216
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_136
timestamp 1719433677
transform 1 0 -233904 0 1 42216
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_137
timestamp 1719433677
transform 1 0 96210 0 1 42616
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_138
timestamp 1719433677
transform 1 0 119666 0 1 42616
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_139
timestamp 1719433677
transform 1 0 137556 0 1 42616
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_140
timestamp 1719433677
transform 0 1 -63730 -1 0 435456
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_141
timestamp 1719433677
transform 0 1 -70394 -1 0 435456
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_142
timestamp 1719433677
transform 0 1 -69882 -1 0 435456
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_143
timestamp 1719433677
transform 0 1 -69370 -1 0 435456
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_144
timestamp 1719433677
transform 0 1 -68858 -1 0 435456
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_145
timestamp 1719433677
transform 0 1 -68346 -1 0 435456
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_146
timestamp 1719433677
transform 0 1 -67834 -1 0 435456
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_147
timestamp 1719433677
transform 0 1 -67322 -1 0 435456
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_148
timestamp 1719433677
transform 0 1 -66810 -1 0 435456
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_149
timestamp 1719433677
transform 0 1 -66298 -1 0 435456
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_150
timestamp 1719433677
transform 0 1 -65786 -1 0 435456
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_151
timestamp 1719433677
transform 0 1 -65274 -1 0 435456
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_152
timestamp 1719433677
transform 0 1 -64762 -1 0 435456
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_153
timestamp 1719433677
transform 0 1 -64250 -1 0 435456
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_154
timestamp 1719433677
transform 0 1 494726 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_155
timestamp 1719433677
transform 0 1 491654 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_156
timestamp 1719433677
transform 0 1 492166 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_157
timestamp 1719433677
transform 0 1 492678 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_158
timestamp 1719433677
transform 0 1 493190 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_159
timestamp 1719433677
transform 0 1 493702 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_160
timestamp 1719433677
transform 0 1 494214 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_161
timestamp 1719433677
transform 0 1 500878 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_162
timestamp 1719433677
transform 0 1 495238 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_163
timestamp 1719433677
transform 0 1 495758 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_164
timestamp 1719433677
transform 0 1 496270 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_165
timestamp 1719433677
transform 0 1 496782 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_166
timestamp 1719433677
transform 0 1 497294 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_167
timestamp 1719433677
transform 0 1 497806 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_168
timestamp 1719433677
transform 0 1 498318 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_169
timestamp 1719433677
transform 0 1 498830 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_170
timestamp 1719433677
transform 0 1 499342 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_171
timestamp 1719433677
transform 0 1 499854 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_172
timestamp 1719433677
transform 0 1 500366 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_173
timestamp 1719433677
transform 0 1 501390 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_174
timestamp 1719433677
transform 0 1 501902 -1 0 435080
box 431918 70502 432946 70630
use cv3_via3_30cut  cv3_via3_30cut_0
timestamp 1719173267
transform 1 0 7000 0 1 3123
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_1
timestamp 1719173267
transform 1 0 6400 0 1 2600
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_2
timestamp 1719173267
transform 1 0 -600 0 1 -75958
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_3
timestamp 1719173267
transform 1 0 5799 0 1 -10237
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_4
timestamp 1719173267
transform 1 0 5201 0 1 -11242
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_5
timestamp 1719173267
transform 1 0 -1200 0 1 -30868
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_6
timestamp 1719173267
transform 1 0 -600 0 1 -31934
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_7
timestamp 1719173267
transform 1 0 599 0 1 -40066
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_8
timestamp 1719173267
transform 1 0 0 0 1 -43270
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_9
timestamp 1719173267
transform 1 0 1200 0 1 -45100
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_10
timestamp 1719173267
transform 1 0 1800 0 1 -47410
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_11
timestamp 1719173267
transform 1 0 2400 0 1 -56536
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_12
timestamp 1719173267
transform 1 0 3000 0 1 -57180
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_13
timestamp 1719173267
transform 1 0 3600 0 1 -58448
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_14
timestamp 1719173267
transform 1 0 4200 0 1 -63972
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_15
timestamp 1719173267
transform 1 0 -2400 0 1 -70442
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_16
timestamp 1719173267
transform 0 1 477954 -1 0 681444
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_17
timestamp 1719173267
transform 0 1 460096 -1 0 680914
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_18
timestamp 1719173267
transform 0 1 413022 -1 0 679672
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_19
timestamp 1719173267
transform 1 0 4356 0 1 -24886
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_20
timestamp 1719173267
transform 0 1 -77428 -1 0 573816
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_21
timestamp 1719173267
transform 0 1 343262 -1 0 679668
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_22
timestamp 1719173267
transform 0 1 319012 -1 0 679672
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_23
timestamp 1719173267
transform 0 1 294998 -1 0 679676
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_24
timestamp 1719173267
transform 0 1 271034 -1 0 679672
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_25
timestamp 1719173267
transform 0 1 364818 -1 0 647802
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_26
timestamp 1719173267
transform 0 1 361570 -1 0 649214
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_27
timestamp 1719173267
transform 0 1 287744 -1 0 649202
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_28
timestamp 1719173267
transform 0 1 286066 -1 0 647624
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_30
timestamp 1719173267
transform 0 1 205274 -1 0 681108
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_31
timestamp 1719173267
transform -1 0 850156 0 -1 205993
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_32
timestamp 1719173267
transform 0 1 173716 -1 0 679678
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_33
timestamp 1719173267
transform 0 1 131634 -1 0 681124
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_34
timestamp 1719173267
transform 0 1 107606 -1 0 680714
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_35
timestamp 1719173267
transform 0 1 83590 -1 0 680310
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_36
timestamp 1719173267
transform 0 1 58436 -1 0 679672
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_37
timestamp 1719173267
transform 0 1 -11574 -1 0 679676
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_38
timestamp 1719173267
transform 0 1 -35220 -1 0 679676
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_39
timestamp 1719173267
transform 0 1 -59256 -1 0 679674
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_40
timestamp 1719173267
transform 0 1 -82954 -1 0 679568
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_41
timestamp 1719173267
transform 0 1 -76934 -1 0 585178
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_42
timestamp 1719173267
transform 0 1 -76938 -1 0 574438
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_43
timestamp 1719173267
transform 0 1 -78452 -1 0 586972
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_44
timestamp 1719173267
transform 0 1 -77946 -1 0 586360
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_45
timestamp 1719173267
transform 0 1 -77424 -1 0 585792
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_46
timestamp 1719173267
transform -1 0 577570 0 -1 125940
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_47
timestamp 1719173267
transform -1 0 579152 0 -1 124678
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_48
timestamp 1719173267
transform -1 0 578620 0 -1 125054
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_49
timestamp 1719173267
transform -1 0 578088 0 -1 125486
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_50
timestamp 1719173267
transform -1 0 575502 0 -1 139940
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_51
timestamp 1719173267
transform -1 0 576020 0 -1 139486
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_52
timestamp 1719173267
transform -1 0 576552 0 -1 139054
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_53
timestamp 1719173267
transform -1 0 577084 0 -1 138678
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_54
timestamp 1719173267
transform -1 0 574484 0 -1 153054
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_55
timestamp 1719173267
transform -1 0 575016 0 -1 152678
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_56
timestamp 1719173267
transform 0 1 -85164 -1 0 643644
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_57
timestamp 1719173267
transform 0 1 -84642 -1 0 643200
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_58
timestamp 1719173267
transform 0 1 -85788 -1 0 656938
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_59
timestamp 1719173267
transform 0 1 -85810 -1 0 656358
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_60
timestamp 1719173267
transform 1 0 -224167 0 1 -82505
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_61
timestamp 1719173267
transform 1 0 -212344 0 1 -79768
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_62
timestamp 1719173267
transform 1 0 -212864 0 1 -80026
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_63
timestamp 1719173267
transform 1 0 -213368 0 1 -80330
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_64
timestamp 1719173267
transform 1 0 -213900 0 1 -80646
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_65
timestamp 1719173267
transform 1 0 -214422 0 1 -80946
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_66
timestamp 1719173267
transform 1 0 -214918 0 1 -81244
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_67
timestamp 1719173267
transform 1 0 -213545 0 1 -72784
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_68
timestamp 1719173267
transform 1 0 -213107 0 1 -75190
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_69
timestamp 1719173267
transform 1 0 -216482 0 1 -80558
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_70
timestamp 1719173267
transform 1 0 -216968 0 1 -80850
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_71
timestamp 1719173267
transform 1 0 -217482 0 1 -81142
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_72
timestamp 1719173267
transform 1 0 -218016 0 1 -81452
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_73
timestamp 1719173267
transform 1 0 -218518 0 1 -81746
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_74
timestamp 1719173267
transform 1 0 -219016 0 1 -82038
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_75
timestamp 1719173267
transform 1 0 -219544 0 1 -82360
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_76
timestamp 1719173267
transform 1 0 -220040 0 1 -82640
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_77
timestamp 1719173267
transform 0 1 -87277 -1 0 582897
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_78
timestamp 1719173267
transform 1 0 1306 0 1 -82348
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_79
timestamp 1719173267
transform 1 0 -462806 0 1 6678
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_80
timestamp 1719173267
transform 1 0 -477170 0 1 6722
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_81
timestamp 1719173267
transform 1 0 -475662 0 1 14499
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_82
timestamp 1719173267
transform 1 0 -463796 0 1 14878
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_83
timestamp 1719173267
transform 1 0 -203501 0 1 -84238
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_84
timestamp 1719173267
transform -1 0 1104171 0 -1 171316
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_85
timestamp 1719173267
transform 0 1 362304 -1 0 585736
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_86
timestamp 1719173267
transform 0 1 360734 -1 0 586234
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_87
timestamp 1719173267
transform 0 1 397228 -1 0 652009
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_88
timestamp 1719173267
transform 0 1 137060 -1 0 644866
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_89
timestamp 1719173267
transform 0 1 134997 -1 0 574460
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_90
timestamp 1719173267
transform 1 0 -220574 0 1 -82958
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_91
timestamp 1719173267
transform 1 0 -75524 0 1 7144
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_92
timestamp 1719173267
transform 1 0 -74040 0 1 15154
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_93
timestamp 1719173267
transform 1 0 -60020 0 1 7144
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_94
timestamp 1719173267
transform 1 0 -60860 0 1 15196
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_95
timestamp 1719173267
transform 0 1 397997 -1 0 644379
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_96
timestamp 1719173267
transform 0 1 414894 -1 0 643171
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_97
timestamp 1719173267
transform 0 1 414540 -1 0 643596
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_98
timestamp 1719173267
transform 0 1 399936 -1 0 643959
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_99
timestamp 1719173267
transform 0 1 324314 -1 0 583451
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_100
timestamp 1719173267
transform 0 -1 454542 1 0 -490434
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_101
timestamp 1719173267
transform 0 -1 454032 1 0 -490054
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_102
timestamp 1719173267
transform 0 -1 453502 1 0 -489628
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_103
timestamp 1719173267
transform 0 -1 453022 1 0 -489226
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_104
timestamp 1719173267
transform 0 -1 446252 1 0 -490440
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_105
timestamp 1719173267
transform 1 0 -214008 0 1 -74447
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_106
timestamp 1719173267
transform 0 1 -82374 -1 0 680186
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_107
timestamp 1719173267
transform 0 1 -58396 -1 0 680572
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_108
timestamp 1719173267
transform 0 -1 451934 1 0 -486020
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_109
timestamp 1719173267
transform 0 -1 451452 1 0 -486414
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_110
timestamp 1719173267
transform 0 -1 450948 1 0 -486816
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_111
timestamp 1719173267
transform 0 -1 450412 1 0 -487218
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_112
timestamp 1719173267
transform 0 -1 449908 1 0 -487636
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_113
timestamp 1719173267
transform 0 -1 449324 1 0 -488024
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_114
timestamp 1719173267
transform 0 -1 448808 1 0 -488414
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_115
timestamp 1719173267
transform 0 -1 448306 1 0 -488836
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_116
timestamp 1719173267
transform 0 -1 447788 1 0 -489206
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_117
timestamp 1719173267
transform 0 -1 447306 1 0 -489600
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_118
timestamp 1719173267
transform 0 -1 446750 1 0 -490016
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_119
timestamp 1719173267
transform 0 1 -34392 -1 0 680972
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_120
timestamp 1719173267
transform 0 -1 181446 1 0 -490452
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_121
timestamp 1719173267
transform 0 1 -10426 -1 0 681352
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_122
timestamp 1719173267
transform 0 1 59610 -1 0 679916
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_123
timestamp 1719173267
transform 0 1 206090 -1 0 680672
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_124
timestamp 1719173267
transform 0 -1 195555 1 0 -489224
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_125
timestamp 1719173267
transform 0 -1 194806 1 0 -489606
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_126
timestamp 1719173267
transform 0 -1 181812 1 0 -490060
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_127
timestamp 1719173267
transform 0 1 471416 -1 0 584342
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_128
timestamp 1719173267
transform 0 1 463578 -1 0 573222
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_129
timestamp 1719173267
transform 0 1 471314 -1 0 575682
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_130
timestamp 1719173267
transform 0 1 470215 -1 0 575178
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_131
timestamp 1719173267
transform 0 1 472856 -1 0 574486
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_132
timestamp 1719173267
transform 0 1 471821 -1 0 575283
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_133
timestamp 1719173267
transform 0 1 472309 -1 0 574909
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_134
timestamp 1719173267
transform 1 0 -409058 0 1 3299
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_135
timestamp 1719173267
transform 1 0 -25814 0 1 -73301
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_136
timestamp 1719173267
transform 0 -1 623304 1 0 -532787
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_137
timestamp 1719173267
transform -1 0 1107800 0 -1 139106
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_138
timestamp 1719173267
transform 1 0 -1800 0 1 -71576
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_139
timestamp 1719173267
transform 1 0 -1200 0 1 -74840
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_140
timestamp 1719173267
transform 1 0 -1800 0 1 -74398
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_141
timestamp 1719173267
transform 1 0 -26365 0 1 -73674
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_142
timestamp 1719173267
transform 1 0 -35326 0 1 -74835
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_143
timestamp 1719173267
transform -1 0 1107239 0 -1 139106
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_144
timestamp 1719173267
transform -1 0 1094602 0 -1 139652
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_145
timestamp 1719173267
transform 1 0 -38505 0 1 -58470
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_146
timestamp 1719173267
transform 1 0 -35961 0 1 -75287
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_147
timestamp 1719173267
transform 1 0 -83366 0 1 -76650
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_148
timestamp 1719173267
transform 1 0 -410233 0 1 529
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_149
timestamp 1719173267
transform 1 0 -409643 0 1 2003
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_150
timestamp 1719173267
transform 0 1 107578 1 0 -476258
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_151
timestamp 1719173267
transform -1 0 764655 0 1 2263
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_152
timestamp 1719173267
transform -1 0 764070 0 1 3559
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_153
timestamp 1719173267
transform 0 1 297660 -1 0 656079
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_154
timestamp 1719173267
transform 1 0 -175373 0 1 2493
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_155
timestamp 1719173267
transform 1 0 -174688 0 1 3789
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_156
timestamp 1719173267
transform 0 1 344004 1 0 -477493
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_157
timestamp 1719173267
transform -1 0 999725 0 1 2523
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_158
timestamp 1719173267
transform -1 0 999240 0 1 3819
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_159
timestamp 1719173267
transform 0 1 108299 -1 0 629624
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_160
timestamp 1719173267
transform 1 0 -179735 0 1 -31549
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_161
timestamp 1719173267
transform 0 1 64455 -1 0 629275
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_162
timestamp 1719173267
transform 1 0 -178346 0 1 -30047
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_163
timestamp 1719173267
transform -1 0 641243 0 -1 166230
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_164
timestamp 1719173267
transform -1 0 652054 0 -1 166307
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_165
timestamp 1719173267
transform -1 0 1093617 0 -1 170922
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_167
timestamp 1719173267
transform 0 1 295107 -1 0 627939
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_168
timestamp 1719173267
transform 0 1 134042 -1 0 577389
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_169
timestamp 1719173267
transform 1 0 -370082 0 1 -80725
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_170
timestamp 1719173267
transform 0 1 105796 -1 0 577390
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_171
timestamp 1719173267
transform 1 0 -340524 0 1 -80716
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_172
timestamp 1719173267
transform 1 0 -399475 0 1 -80857
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_173
timestamp 1719173267
transform 0 1 75051 -1 0 577254
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_174
timestamp 1719173267
transform 0 1 46845 -1 0 577255
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_175
timestamp 1719173267
transform 1 0 -429034 0 1 -80855
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_176
timestamp 1719173267
transform 0 1 134635 -1 0 573831
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_177
timestamp 1719173267
transform -1 0 796858 0 -1 100611
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_178
timestamp 1719173267
transform 0 1 471788 -1 0 584816
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_179
timestamp 1719173267
transform 0 1 104893 -1 0 574445
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_180
timestamp 1719173267
transform 0 1 105242 -1 0 573821
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_181
timestamp 1719173267
transform 0 1 45904 -1 0 574442
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_182
timestamp 1719173267
transform 0 1 76043 -1 0 574438
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_183
timestamp 1719173267
transform 0 1 75669 -1 0 573809
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_184
timestamp 1719173267
transform 0 1 46273 -1 0 573813
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_185
timestamp 1719173267
transform 0 1 14805 -1 0 573191
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_186
timestamp 1719173267
transform 0 1 16904 -1 0 572579
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_187
timestamp 1719173267
transform 0 1 15218 -1 0 584953
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_188
timestamp 1719173267
transform 0 1 16516 -1 0 602592
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_189
timestamp 1719173267
transform 0 1 -86696 -1 0 578212
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_190
timestamp 1719173267
transform -1 0 571436 0 -1 154669
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_191
timestamp 1719173267
transform 0 1 297690 -1 0 586716
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_192
timestamp 1719173267
transform 0 1 435382 -1 0 574530
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_193
timestamp 1719173267
transform 1 0 -105458 0 1 -73822
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_194
timestamp 1719173267
transform 0 1 324219 -1 0 584061
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_195
timestamp 1719173267
transform 0 1 295064 -1 0 585403
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_196
timestamp 1719173267
transform 1 0 -179722 0 1 -71716
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_197
timestamp 1719173267
transform 0 1 296544 -1 0 587128
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_198
timestamp 1719173267
transform 1 0 -131273 0 1 -48378
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_199
timestamp 1719173267
transform 0 1 344286 -1 0 585928
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_200
timestamp 1719173267
transform 0 1 339684 -1 0 587596
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_201
timestamp 1719173267
transform 0 1 296131 -1 0 628285
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_202
timestamp 1719173267
transform 1 0 -178978 0 1 -70034
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_203
timestamp 1719173267
transform 0 1 455476 -1 0 572580
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_204
timestamp 1719173267
transform 0 1 463566 -1 0 587104
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_205
timestamp 1719173267
transform 0 1 455542 -1 0 587076
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_206
timestamp 1719173267
transform 0 1 436467 -1 0 575985
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_207
timestamp 1719173267
transform -1 0 1094026 0 -1 126270
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_208
timestamp 1719173267
transform 1 0 -40104 0 1 -70934
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_209
timestamp 1719173267
transform 1 0 -82926 0 1 -75189
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_210
timestamp 1719173267
transform 1 0 -82564 0 1 -73992
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_211
timestamp 1719173267
transform 1 0 -534424 0 1 -2800
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_212
timestamp 1719173267
transform 1 0 -534002 0 1 -2392
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_213
timestamp 1719173267
transform 1 0 -535224 0 1 -14992
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_214
timestamp 1719173267
transform 1 0 -534826 0 1 -13848
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_215
timestamp 1719173267
transform 1 0 -531590 0 1 -30160
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_216
timestamp 1719173267
transform 1 0 -531984 0 1 -31094
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_217
timestamp 1719173267
transform 1 0 -532398 0 1 -41446
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_218
timestamp 1719173267
transform 1 0 -532802 0 1 -42600
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_219
timestamp 1719173267
transform 1 0 -533204 0 1 -43948
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_220
timestamp 1719173267
transform 1 0 -533588 0 1 -44898
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_221
timestamp 1719173267
transform 1 0 -533992 0 1 -55464
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_222
timestamp 1719173267
transform 1 0 -534406 0 1 -56614
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_223
timestamp 1719173267
transform 1 0 -534784 0 1 -57944
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_224
timestamp 1719173267
transform 1 0 -535204 0 1 -59016
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_225
timestamp 1719173267
transform 0 1 63606 -1 0 657086
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_226
timestamp 1719173267
transform 0 1 64308 -1 0 655584
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_227
timestamp 1719173267
transform -1 0 765245 0 1 789
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_228
timestamp 1719173267
transform 0 1 108544 1 0 -477796
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_229
timestamp 1719173267
transform 1 0 -175863 0 1 1019
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_230
timestamp 1719173267
transform 0 1 298508 -1 0 657623
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_231
timestamp 1719173267
transform -1 0 1000515 0 1 1049
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_232
timestamp 1719173267
transform 0 1 342967 1 0 -475961
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_233
timestamp 1719173267
transform 0 1 198008 -1 0 679678
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_234
timestamp 1719173267
transform -1 0 852592 0 -1 205116
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_235
timestamp 1719173267
transform -1 0 851772 0 -1 205535
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_236
timestamp 1719173267
transform -1 0 850970 0 -1 206006
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_237
timestamp 1719173267
transform -1 0 851778 0 -1 142811
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_238
timestamp 1719173267
transform -1 0 850930 0 -1 199373
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_239
timestamp 1719173267
transform -1 0 850974 0 -1 195950
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_240
timestamp 1719173267
transform -1 0 852608 0 -1 187916
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_241
timestamp 1719173267
transform -1 0 850130 0 -1 183276
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_242
timestamp 1719173267
transform -1 0 850130 0 -1 179798
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_243
timestamp 1719173267
transform -1 0 851804 0 -1 171875
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_244
timestamp 1719173267
transform -1 0 850135 0 -1 151967
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_245
timestamp 1719173267
transform -1 0 850968 0 -1 147264
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_246
timestamp 1719173267
transform -1 0 850153 0 -1 111268
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_247
timestamp 1719173267
transform -1 0 852586 0 -1 138217
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_248
timestamp 1719173267
transform -1 0 850967 0 -1 124219
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_249
timestamp 1719173267
transform -1 0 1093513 0 -1 153156
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_250
timestamp 1719173267
transform -1 0 1094062 0 -1 152618
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_251
timestamp 1719173267
transform -1 0 1094588 0 -1 152130
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_252
timestamp 1719173267
transform -1 0 1097645 0 -1 138574
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_253
timestamp 1719173267
transform 0 1 207056 -1 0 679670
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_254
timestamp 1719173267
transform 0 1 197058 -1 0 681512
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_255
timestamp 1719173267
transform 0 1 174616 -1 0 681528
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_256
timestamp 1719173267
transform 0 1 270064 -1 0 681428
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_257
timestamp 1719173267
transform 0 1 294064 -1 0 680948
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_258
timestamp 1719173267
transform 0 1 318090 -1 0 680558
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_259
timestamp 1719173267
transform 0 1 342102 -1 0 680134
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_260
timestamp 1719173267
transform 0 1 412070 -1 0 681208
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_261
timestamp 1719173267
transform 0 1 436064 -1 0 681474
box 566656 91154 566956 91980
use cv3_via4_2cut  cv3_via4_2cut_0
timestamp 1717863568
transform 0 1 571823 -1 0 16443
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_1
timestamp 1717863568
transform 0 1 572674 -1 0 12880
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_2
timestamp 1717863568
transform 0 1 572430 -1 0 34846
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_3
timestamp 1717863568
transform 0 1 570978 -1 0 75518
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_4
timestamp 1717863568
transform 1 0 6070 0 1 29202
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_5
timestamp 1717863568
transform 1 0 5542 0 1 50214
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_6
timestamp 1717863568
transform 1 0 7316 0 1 72198
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_7
timestamp 1717863568
transform 1 0 7308 0 1 93208
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_8
timestamp 1717863568
transform 0 1 573630 -1 0 76839
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_9
timestamp 1717863568
transform 0 1 573021 -1 0 55840
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_10
timestamp 1717863568
transform 0 1 570966 -1 0 54890
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_11
timestamp 1717863568
transform 1 0 4930 0 1 92192
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_12
timestamp 1717863568
transform 1 0 4910 0 1 71200
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_13
timestamp 1717863568
transform 0 1 6958 -1 0 30910
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_14
timestamp 1717863568
transform 0 1 6958 -1 0 51912
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_15
timestamp 1717863568
transform 0 1 570972 -1 0 33892
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_16
timestamp 1717863568
transform 0 1 572680 -1 0 33528
box 0 0 688 368
use cv3_via_3cut  cv3_via_3cut_0
timestamp 1719452912
transform 1 0 1108 0 1 1311
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_1
timestamp 1719452912
transform 1 0 0 0 1 1900
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_2
timestamp 1719452912
transform 1 0 102 0 1 1824
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_3
timestamp 1719452912
transform 1 0 215 0 1 1751
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_4
timestamp 1719452912
transform 1 0 329 0 1 1674
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_5
timestamp 1719452912
transform 1 0 439 0 1 1600
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_6
timestamp 1719452912
transform 1 0 546 0 1 1533
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_7
timestamp 1719452912
transform 1 0 664 0 1 1463
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_8
timestamp 1719452912
transform 1 0 766 0 1 1394
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_9
timestamp 1719452912
transform 1 0 552403 0 1 -48894
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_10
timestamp 1719452912
transform 1 0 554081 0 1 -50692
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_11
timestamp 1719452912
transform 1 0 1216 0 1 1242
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_12
timestamp 1719452912
transform 1 0 1893 0 1 802
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_13
timestamp 1719452912
transform 1 0 1332 0 1 1164
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_14
timestamp 1719452912
transform 1 0 1438 0 1 1098
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_15
timestamp 1719452912
transform 1 0 1560 0 1 1027
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_16
timestamp 1719452912
transform 1 0 1674 0 1 953
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_17
timestamp 1719452912
transform 1 0 1783 0 1 876
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_18
timestamp 1719452912
transform 1 0 553969 0 1 -50568
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_19
timestamp 1719452912
transform 1 0 553861 0 1 -50452
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_20
timestamp 1719452912
transform 1 0 553753 0 1 -50334
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_21
timestamp 1719452912
transform 1 0 553635 0 1 -50214
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_22
timestamp 1719452912
transform 1 0 553519 0 1 -50094
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_23
timestamp 1719452912
transform 1 0 553407 0 1 -49980
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_24
timestamp 1719452912
transform 1 0 553297 0 1 -49864
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_25
timestamp 1719452912
transform 1 0 553185 0 1 -49756
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_26
timestamp 1719452912
transform 1 0 553071 0 1 -49628
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_27
timestamp 1719452912
transform 1 0 552963 0 1 -49516
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_28
timestamp 1719452912
transform 1 0 552845 0 1 -49392
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_29
timestamp 1719452912
transform 1 0 552725 0 1 -49246
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_30
timestamp 1719452912
transform 1 0 552625 0 1 -49144
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_31
timestamp 1719452912
transform 1 0 552515 0 1 -49026
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_32
timestamp 1719452912
transform 1 0 557475 0 1 -49144
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_33
timestamp 1719452912
transform 1 0 557117 0 1 -48774
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_34
timestamp 1719452912
transform 1 0 557237 0 1 -48894
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_35
timestamp 1719452912
transform 1 0 557355 0 1 -49012
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_36
timestamp 1719452912
transform 1 0 558915 0 1 -50572
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_37
timestamp 1719452912
transform 1 0 557599 0 1 -49258
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_38
timestamp 1719452912
transform 1 0 557717 0 1 -49372
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_39
timestamp 1719452912
transform 1 0 557833 0 1 -49488
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_40
timestamp 1719452912
transform 1 0 557961 0 1 -49606
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_41
timestamp 1719452912
transform 1 0 558081 0 1 -49726
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_42
timestamp 1719452912
transform 1 0 558193 0 1 -49846
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_43
timestamp 1719452912
transform 1 0 558317 0 1 -49968
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_44
timestamp 1719452912
transform 1 0 558441 0 1 -50092
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_45
timestamp 1719452912
transform 1 0 558549 0 1 -50210
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_46
timestamp 1719452912
transform 1 0 558679 0 1 -50326
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_47
timestamp 1719452912
transform 1 0 558793 0 1 -50454
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_48
timestamp 1719452912
transform 1 0 559473 0 1 3758
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_49
timestamp 1719452912
transform 1 0 559111 0 1 3408
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_50
timestamp 1719452912
transform 1 0 559235 0 1 3534
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_51
timestamp 1719452912
transform 1 0 559353 0 1 3638
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_52
timestamp 1719452912
transform 1 0 560793 0 1 5078
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_53
timestamp 1719452912
transform 1 0 559593 0 1 3878
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_54
timestamp 1719452912
transform 1 0 559713 0 1 3998
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_55
timestamp 1719452912
transform 1 0 559833 0 1 4118
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_56
timestamp 1719452912
transform 1 0 559953 0 1 4238
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_57
timestamp 1719452912
transform 1 0 560073 0 1 4358
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_58
timestamp 1719452912
transform 1 0 560193 0 1 4478
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_59
timestamp 1719452912
transform 1 0 560313 0 1 4598
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_60
timestamp 1719452912
transform 1 0 560433 0 1 4718
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_61
timestamp 1719452912
transform 1 0 560553 0 1 4838
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_62
timestamp 1719452912
transform 1 0 560673 0 1 4958
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_63
timestamp 1719452912
transform 1 0 560913 0 1 5198
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_64
timestamp 1719452912
transform 0 1 440340 -1 0 70673
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_65
timestamp 1719452912
transform 0 1 440118 -1 0 71029
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_66
timestamp 1719452912
transform 0 1 440184 -1 0 70909
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_67
timestamp 1719452912
transform 0 1 440262 -1 0 70787
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_68
timestamp 1719452912
transform 0 1 445504 -1 0 70381
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_69
timestamp 1719452912
transform 0 1 445726 -1 0 70693
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_70
timestamp 1719452912
transform 0 1 445650 -1 0 70577
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_71
timestamp 1719452912
transform 0 1 445578 -1 0 70481
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_72
timestamp 1719452912
transform 0 1 450136 -1 0 70787
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_73
timestamp 1719452912
transform 0 1 450356 -1 0 71109
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_74
timestamp 1719452912
transform 0 1 450284 -1 0 70995
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_75
timestamp 1719452912
transform 0 1 450214 -1 0 70883
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_76
timestamp 1719452912
transform 0 1 454749 -1 0 71111
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_77
timestamp 1719452912
transform 0 1 454526 -1 0 70754
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_78
timestamp 1719452912
transform 0 1 454604 -1 0 70847
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_80
timestamp 1719452912
transform 1 0 534711 0 1 -95842
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_81
timestamp 1719452912
transform 1 0 532921 0 1 -96578
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_82
timestamp 1719452912
transform 1 0 533025 0 1 -96502
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_83
timestamp 1719452912
transform 1 0 533143 0 1 -96430
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_84
timestamp 1719452912
transform 1 0 533255 0 1 -96362
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_85
timestamp 1719452912
transform 1 0 533703 0 1 -96286
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_86
timestamp 1719452912
transform 1 0 533815 0 1 -96214
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_87
timestamp 1719452912
transform 1 0 533925 0 1 -96136
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_88
timestamp 1719452912
transform 1 0 534379 0 1 -96060
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_89
timestamp 1719452912
transform 1 0 534489 0 1 -95988
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_90
timestamp 1719452912
transform 1 0 534599 0 1 -95916
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_91
timestamp 1719452912
transform 1 0 535721 0 1 -95474
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_92
timestamp 1719452912
transform 1 0 535159 0 1 -95770
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_93
timestamp 1719452912
transform 1 0 535269 0 1 -95692
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_94
timestamp 1719452912
transform 1 0 535381 0 1 -95618
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_95
timestamp 1719452912
transform 1 0 535607 0 1 -95546
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_96
timestamp 1719452912
transform 1 0 536379 0 1 -95172
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_97
timestamp 1719452912
transform 1 0 536165 0 1 -95250
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_98
timestamp 1719452912
transform 1 0 535941 0 1 -95402
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_99
timestamp 1719452912
transform 1 0 536051 0 1 -95326
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_100
timestamp 1719452912
transform 1 0 536607 0 1 -95030
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_101
timestamp 1719452912
transform 1 0 536499 0 1 -95106
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_102
timestamp 1719452912
transform 1 0 538183 0 1 -94214
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_103
timestamp 1719452912
transform 1 0 536837 0 1 -94956
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_104
timestamp 1719452912
transform 1 0 536951 0 1 -94882
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_105
timestamp 1719452912
transform 1 0 537173 0 1 -94806
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_106
timestamp 1719452912
transform 1 0 537281 0 1 -94736
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_107
timestamp 1719452912
transform 1 0 537397 0 1 -94658
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_108
timestamp 1719452912
transform 1 0 537619 0 1 -94586
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_109
timestamp 1719452912
transform 1 0 537729 0 1 -94512
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_110
timestamp 1719452912
transform 1 0 537845 0 1 -94438
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_111
timestamp 1719452912
transform 1 0 537961 0 1 -94362
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_112
timestamp 1719452912
transform 1 0 538067 0 1 -94288
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_113
timestamp 1719452912
transform 1 0 538629 0 1 -93920
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_114
timestamp 1719452912
transform 1 0 538293 0 1 -94138
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_115
timestamp 1719452912
transform 1 0 538405 0 1 -94066
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_116
timestamp 1719452912
transform 1 0 538519 0 1 -93994
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_117
timestamp 1719452912
transform 1 0 540979 0 1 -93472
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_118
timestamp 1719452912
transform 1 0 539749 0 1 -93842
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_119
timestamp 1719452912
transform 1 0 539861 0 1 -93772
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_120
timestamp 1719452912
transform 1 0 539973 0 1 -93698
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_121
timestamp 1719452912
transform 1 0 540755 0 1 -93620
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_122
timestamp 1719452912
transform 1 0 540867 0 1 -93550
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_123
timestamp 1719452912
transform 1 0 543221 0 1 -93106
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_124
timestamp 1719452912
transform 1 0 542103 0 1 -93398
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_125
timestamp 1719452912
transform 1 0 542215 0 1 -93328
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_126
timestamp 1719452912
transform 1 0 542997 0 1 -93252
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_127
timestamp 1719452912
transform 1 0 543109 0 1 -93180
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_128
timestamp 1719452912
transform 1 0 544789 0 1 -92736
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_129
timestamp 1719452912
transform 1 0 544123 0 1 -93030
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_130
timestamp 1719452912
transform 1 0 544227 0 1 -92958
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_131
timestamp 1719452912
transform 1 0 544569 0 1 -92882
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_132
timestamp 1719452912
transform 1 0 544675 0 1 -92812
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_133
timestamp 1719452912
transform 1 0 164123 0 1 -105170
box 10601 106968 10663 107172
use cv3_via_3cut  cv3_via_3cut_134
timestamp 1719452912
transform 1 0 221684 0 1 -104901
box 10601 106968 10663 107172
use cv3_via_30cut  cv3_via_30cut_0
timestamp 1719247715
transform 1 0 478530 0 1 -93394
box 14334 104924 14594 105610
use cv3_via_30cut  cv3_via_30cut_10
timestamp 1719247715
transform 1 0 349699 0 1 -46536
box 14334 104924 14594 105610
use cv3_via_30cut  cv3_via_30cut_11
timestamp 1719247715
transform 1 0 350246 0 1 -46181
box 14334 104924 14594 105610
use cv3_via_30cut  cv3_via_30cut_12
timestamp 1719247715
transform 1 0 391188 0 1 -44926
box 14334 104924 14594 105610
use cv3_via_30cut  cv3_via_30cut_13
timestamp 1719247715
transform 1 0 391849 0 1 -44917
box 14334 104924 14594 105610
use cv3_via_30cut  cv3_via_30cut_14
timestamp 1719247715
transform 1 0 391520 0 1 -44919
box 14334 104924 14594 105610
use cv3_via_30cut  cv3_via_30cut_15
timestamp 1719247715
transform 1 0 172426 0 1 -51563
box 14334 104924 14594 105610
use cv3_via_30cut  cv3_via_30cut_16
timestamp 1719247715
transform 1 0 172435 0 1 -47133
box 14334 104924 14594 105610
use cv3_via_30cut  cv3_via_30cut_17
timestamp 1719247715
transform 1 0 171666 0 1 -50563
box 14334 104924 14594 105610
use simple_analog_mux_sel1v8  simple_analog_mux_sel1v8_0 ../dependencies/sky130_ef_ip__analog_switches/mag
timestamp 1724439832
transform 1 0 187386 0 -1 56125
box -46 -2540 3538 3648
use simple_analog_mux_sel1v8  simple_analog_mux_sel1v8_1
timestamp 1724439832
transform -1 0 421022 0 -1 49627
box -46 -2540 3538 3648
use simple_switch_array_3  simple_switch_array_3_0
timestamp 1724444265
transform 1 0 143682 0 1 77405
box -186 881 12599 5129
use simple_switch_array_3  simple_switch_array_3_1
timestamp 1724444265
transform 1 0 199244 0 1 77541
box -186 881 12599 5129
use simple_switch_array_3  simple_switch_array_3_2
timestamp 1724444265
transform 1 0 376428 0 1 77535
box -186 881 12599 5129
use simple_switch_array_3  simple_switch_array_3_3
timestamp 1724444265
transform 1 0 436018 0 1 77601
box -186 881 12599 5129
use simple_switch_array_6  simple_switch_array_6_0
timestamp 1724444338
transform 1 0 215584 0 1 77523
box -664 858 29188 5129
use simple_switch_array_8  simple_switch_array_8_0
timestamp 1724444186
transform 1 0 454460 0 1 77703
box -974 857 40892 5129
use simple_switch_array_15  simple_switch_array_15_0
timestamp 1726771202
transform 0 1 338541 -1 0 44143
box -12973 3053 29596 13997
use simple_switch_array_16  simple_switch_array_16_0
timestamp 1731205139
transform 1 0 548258 0 1 61913
box -412 -1454 19634 19103
use simple_switch_array_32  simple_switch_array_32_0
timestamp 1724447141
transform -1 0 281616 0 -1 62050
box -935 397 44410 19364
use simple_switch_array_53  simple_switch_array_53_0
timestamp 1724444698
transform 1 0 366085 0 1 61911
box -843 412 140525 16287
use sky130_ajc_ip__brownout  sky130_ajc_ip__brownout_0 ../dependencies/sky130_ajc_ip__brownout/mag
timestamp 1713419710
transform 1 0 37628 0 1 15381
box -1604 -1987 43293 41283
use sky130_ak_ip__cmos_vref  sky130_ak_ip__cmos_vref_0 ../dependencies/sky130_ak_ip__cmos_vref/mag
timestamp 1721067183
transform 0 -1 395482 1 0 37455
box 8587 -19903 21921 206
use sky130_ak_ip__comparator  sky130_ak_ip__comparator_0 ../dependencies/sky130_ak_ip__comparator/mag
timestamp 1738083055
transform 0 1 326450 -1 0 57962
box -1900 -33700 39700 13700
use sky130_am_ip__ldo_01v8  sky130_am_ip__ldo_01v8_0 ../dependencies/sky130_am_ip__ldo_01v8/mag
timestamp 1721052427
transform 0 1 378665 -1 0 48529
box 4253 -10775 28439 6899
use sky130_cw_ip__bandgap_nobias  sky130_cw_ip__bandgap_nobias_0 ../dependencies/sky130_cw_ip/mag
timestamp 1731269207
transform -1 0 474518 0 1 44954
box -396 12 42048 14837
use sky130_ef_ip__biasgen4  sky130_ef_ip__biasgen4_0 ../dependencies/sky130_ef_ip__biasgen/mag
timestamp 1732763842
transform 1 0 363572 0 1 7300
box -67 -505 119540 10896
use sky130_ef_ip__cdac3v_12bit  sky130_ef_ip__cdac3v_12bit_0 ../dependencies/sky130_ef_ip__cdac3v_12bit/mag
timestamp 1731117925
transform 1 0 81345 0 -1 23588
box 52849 -36568 89580 15691
use sky130_ef_ip__cdac3v_12bit  sky130_ef_ip__cdac3v_12bit_1
timestamp 1731117925
transform 1 0 140297 0 -1 23726
box 52849 -36568 89580 15691
use sky130_ef_ip__idac3v_8bit  sky130_ef_ip__idac3v_8bit_0 ../dependencies/sky130_ef_ip__biasgen/mag
timestamp 1724460830
transform 0 1 485688 1 0 11088
box -1186 -1691 49914 35112
use sky130_ef_ip__rdac3v_8bit  sky130_ef_ip__rdac3v_8bit_0 ../dependencies/sky130_ef_ip__rdac3v_8bit/mag
timestamp 1718228761
transform 0 1 109414 1 0 11128
box -200 -200 25939 21270
use sky130_ef_ip__rdac3v_8bit  sky130_ef_ip__rdac3v_8bit_1
timestamp 1718228761
transform 0 -1 105610 1 0 11128
box -200 -200 25939 21270
use sky130_ef_ip__rheostat_8bit  sky130_ef_ip__rheostat_8bit_0 ../dependencies/sky130_ef_ip__rheostat_8bit/mag
timestamp 1716082924
transform 0 1 179122 1 0 81272
box -200 -4 25939 16904
use sky130_ef_ip__rheostat_8bit  sky130_ef_ip__rheostat_8bit_2
timestamp 1716082924
transform 0 1 413200 1 0 80778
box -200 -4 25939 16904
use sky130_ef_ip__rheostat_8bit  sky130_ef_ip__rheostat_8bit_3
timestamp 1716082924
transform 0 -1 409876 1 0 80838
box -200 -4 25939 16904
use sky130_ef_ip__rheostat_8bit  sky130_ef_ip__rheostat_8bit_4
timestamp 1716082924
transform 0 -1 175498 1 0 81290
box -200 -4 25939 16904
use sky130_ef_ip__scomp3v  sky130_ef_ip__scomp3v_0 ../dependencies/sky130_ef_ip__ccomp3v/mag
timestamp 1731034391
transform -1 0 186430 0 -1 32072
box -58 -3122 11186 4094
use sky130_ef_ip__scomp3v  sky130_ef_ip__scomp3v_1
timestamp 1731034391
transform -1 0 243850 0 -1 32240
box -58 -3122 11186 4094
use sky130_fd_io__top_pwrdetv2  sky130_fd_io__top_pwrdetv2_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1733158100
transform 0 1 86014 -1 0 60724
box 282 0 10856 40000
use sky130_fd_io__top_pwrdetv2  sky130_fd_io__top_pwrdetv2_1
timestamp 1733158100
transform 0 1 86014 -1 0 48806
box 282 0 10856 40000
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_0
array 0 0 -2720 0 9 2579
timestamp 1721093827
transform 0 1 320837 1 0 61339
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_1
array 0 2 -3766 0 5 -2724
timestamp 1721093827
transform -1 0 374783 0 -1 23167
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_2
array 0 0 2732 0 15 2564
timestamp 1721093827
transform 0 1 298069 1 0 11908
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_3
array 0 0 -2720 0 9 2579
timestamp 1721093827
transform 0 1 320736 1 0 67370
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_4
array 0 0 2746 0 14 2533
timestamp 1721093827
transform 0 1 43830 1 0 59986
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_5
array 0 0 -2720 0 9 2579
timestamp 1721093827
transform 0 1 294450 1 0 67310
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_6
array 0 0 -2720 0 9 2579
timestamp 1721093827
transform 0 1 321913 1 0 77136
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_7
array 0 0 -2720 0 9 2579
timestamp 1721093827
transform 0 1 294487 1 0 61339
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_8
array 0 0 2732 0 15 2564
timestamp 1721093827
transform 0 1 297993 -1 0 14956
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_9
array 0 1 3268 0 4 2588
timestamp 1721093827
transform 0 1 417124 -1 0 57339
box -1349 -1081 1371 1081
use sky130_icrg_ip__ulpcomp2  sky130_icrg_ip__ulpcomp2_0 ../dependencies/sky130_icrg_ip__ulpcomp/mag
timestamp 1720377809
transform 0 1 372127 -1 0 57532
box -625 -8056 8504 1566
use sky130_iic_ip__audiodac_drv_lite  sky130_iic_ip__audiodac_drv_lite_0 ../dependencies/sky130_iic_ip__audiodac_lite/mag
timestamp 1731463845
transform 1 0 257286 0 1 11406
box -316 -300 9632 28678
use sky130_od_ip__tempsensor_ext_vp  sky130_od_ip__tempsensor_ext_vp_0 ../dependencies/sky130_od_ip__tempsensor/mag
timestamp 1724531563
transform -1 0 185196 0 1 57134
box -584 -5030 6610 3202
use sky130_pa_ip__instramp  sky130_pa_ip__instramp_0 ../dependencies/sky130_pa_ip__instramp/mag
timestamp 1731773078
transform 0 -1 88658 1 0 78128
box 0 0 29566 40042
use sky130_pa_ip__instramp  sky130_pa_ip__instramp_1
timestamp 1731773078
transform 0 -1 550776 1 0 80884
box 0 0 29566 40042
use sky130_sw_ip__por  sky130_sw_ip__por_0 ../dependencies/sky130_sw_ip__por/mag
timestamp 1731723950
transform 1 0 390789 0 1 321922
box 2366 -300396 39669 -277894
use sky130_td_ip__opamp_hp_narrow  sky130_td_ip__opamp_hp_narrow_0 ../dependencies/sky130_td_ip__opamp_hp/mag
timestamp 1731177145
transform 1 0 207046 0 -1 100322
box -7724 -6929 43180 16206
use sky130_td_ip__opamp_hp_narrow  sky130_td_ip__opamp_hp_narrow_1
timestamp 1731177145
transform -1 0 147908 0 -1 100076
box -7724 -6929 43180 16206
use sky130_td_ip__opamp_hp_narrow  sky130_td_ip__opamp_hp_narrow_2
timestamp 1731177145
transform -1 0 382230 0 -1 100570
box -7724 -6929 43180 16206
use sky130_td_ip__opamp_hp_narrow  sky130_td_ip__opamp_hp_narrow_3
timestamp 1731177145
transform 1 0 442290 0 -1 100618
box -7724 -6929 43180 16206
use sky130_vbl_ip__overvoltage  sky130_vbl_ip__overvoltage_0 ../dependencies/sky130_vbl_ip__overvoltage/mag
timestamp 1714660490
transform 1 0 454156 0 1 25528
box -18218 -4002 24405 17489
use switch_array_2  switch_array_2_0
timestamp 1724444975
transform 1 0 274190 0 -1 30916
box -328 -1310 7820 11108
use switch_array_2  switch_array_2_1
timestamp 1724444975
transform 1 0 532088 0 1 22356
box -328 -1310 7820 11108
use switch_array_2  switch_array_2_2
timestamp 1724444975
transform 1 0 532117 0 1 35921
box -328 -1310 7820 11108
use switch_array_2  switch_array_2_3
timestamp 1724444975
transform 0 1 530679 -1 0 58404
box -328 -1310 7820 11108
use switch_array_4  switch_array_4_0
timestamp 1724443940
transform 0 1 91578 1 0 91436
box -328 -1318 15746 11108
use switch_array_4  switch_array_4_1
timestamp 1724443940
transform 0 1 267480 1 0 92050
box -328 -1318 15746 11108
use switch_array_4  switch_array_4_2
timestamp 1724443940
transform 0 1 316082 1 0 91798
box -328 -1318 15746 11108
use switch_array_4  switch_array_4_3
timestamp 1724443940
transform 0 -1 504312 1 0 91760
box -328 -1318 15746 11108
use switch_array_4  switch_array_4_4
timestamp 1724443940
transform 1 0 543936 0 1 22362
box -328 -1318 15746 11108
use switch_array_4  switch_array_4_5
timestamp 1724443940
transform 1 0 544236 0 1 35749
box -328 -1318 15746 11108
use switch_array_4  switch_array_4_6
timestamp 1724443940
transform 1 0 13050 0 1 78416
box -328 -1318 15746 11108
use switch_array_4  switch_array_4_7
timestamp 1724443940
transform 1 0 13206 0 1 22025
box -328 -1318 15746 11108
use switch_array_4  switch_array_4_8
timestamp 1724443940
transform 1 0 552936 0 1 83303
box -328 -1318 15746 11108
use switch_array_4  switch_array_4_9
timestamp 1724443940
transform 1 0 545086 0 1 48986
box -328 -1318 15746 11108
use switch_array_4  switch_array_4_10
timestamp 1724443940
transform 1 0 13206 0 1 50217
box -328 -1318 15746 11108
use switch_array_4  switch_array_4_11
timestamp 1724443940
transform 1 0 13206 0 1 36221
box -328 -1318 15746 11108
use switch_array_14  switch_array_14_1
timestamp 1724444054
transform 0 -1 311182 1 0 77138
box -405 0 31801 23215
use switch_array_18  switch_array_18_0
timestamp 1720191374
transform 1 0 14838 0 1 90894
box -351 -1000 28728 17274
<< labels >>
flabel metal4 368 0 496 300 0 FreeSans 240 90 0 0 gpio5_4
port 1 nsew
flabel metal4 880 0 1008 300 0 FreeSans 240 90 0 0 gpio5_5
port 2 nsew
flabel metal4 1392 0 1520 300 0 FreeSans 240 90 0 0 gpio5_6
port 3 nsew
flabel metal4 1904 0 2032 300 0 FreeSans 240 90 0 0 gpio5_7
port 4 nsew
flabel metal4 2416 0 2544 300 0 FreeSans 240 90 0 0 gpio6_0
port 5 nsew
flabel metal4 3440 0 3568 300 0 FreeSans 240 90 0 0 gpio6_2
port 7 nsew
flabel metal4 3952 0 4080 300 0 FreeSans 240 90 0 0 gpio6_3
port 8 nsew
flabel metal4 4464 0 4592 300 0 FreeSans 240 90 0 0 left_vref
port 9 nsew
flabel metal4 4976 0 5104 300 0 FreeSans 240 90 0 0 gpio6_4
port 10 nsew
flabel metal4 5488 0 5616 300 0 FreeSans 240 90 0 0 gpio6_5
port 11 nsew
flabel metal4 6000 0 6128 300 0 FreeSans 240 90 0 0 gpio6_6
port 12 nsew
flabel metal4 6512 0 6640 300 0 FreeSans 240 90 0 0 gpio6_7
port 13 nsew
flabel metal2 7024 0 7052 300 0 FreeSans 240 90 0 0 adc_refl_to_gpio6_7[1]
port 14 nsew
flabel metal2 7136 0 7164 300 0 FreeSans 240 90 0 0 adc_refl_to_gpio6_7[0]
port 15 nsew
flabel metal2 7248 0 7276 300 0 FreeSans 240 90 0 0 adc_refh_to_gpio6_6[1]
port 16 nsew
flabel metal2 7360 0 7388 300 0 FreeSans 240 90 0 0 adc_refh_to_gpio6_6[0]
port 17 nsew
flabel metal2 7472 0 7500 300 0 FreeSans 240 90 0 0 adc1_to_gpio6_5[1]
port 18 nsew
flabel metal2 7584 0 7612 300 0 FreeSans 240 90 0 0 adc1_to_gpio6_5[0]
port 19 nsew
flabel metal2 7696 0 7724 300 0 FreeSans 240 90 0 0 adc0_to_gpio6_4[1]
port 20 nsew
flabel metal2 7808 0 7836 300 0 FreeSans 240 90 0 0 adc0_to_gpio6_4[0]
port 21 nsew
flabel metal2 7920 0 7948 300 0 FreeSans 240 90 0 0 comp_p_to_gpio6_2[1]
port 22 nsew
flabel metal2 8032 0 8060 300 0 FreeSans 240 90 0 0 comp_p_to_gpio6_2[0]
port 23 nsew
flabel metal2 8144 0 8172 300 0 FreeSans 240 90 0 0 comp_n_to_gpio6_3[1]
port 24 nsew
flabel metal2 8256 0 8284 300 0 FreeSans 240 90 0 0 comp_n_to_gpio6_3[0]
port 25 nsew
flabel metal2 8368 0 8396 300 0 FreeSans 240 90 0 0 ulpcomp_n_to_gpio6_1[1]
port 26 nsew
flabel metal2 8480 0 8508 300 0 FreeSans 240 90 0 0 ulpcomp_n_to_gpio6_1[0]
port 27 nsew
flabel metal2 8592 0 8620 300 0 FreeSans 240 90 0 0 ulpcomp_p_to_gpio6_0[1]
port 28 nsew
flabel metal2 8704 0 8732 300 0 FreeSans 240 90 0 0 ulpcomp_p_to_gpio6_0[0]
port 29 nsew
flabel metal2 8816 0 8844 300 0 FreeSans 240 90 0 0 left_instramp_n_to_gpio5_7[1]
port 30 nsew
flabel metal2 8928 0 8956 300 0 FreeSans 240 90 0 0 left_instramp_n_to_gpio5_7[0]
port 31 nsew
flabel metal2 9040 0 9068 300 0 FreeSans 240 90 0 0 left_instramp_p_to_gpio5_6[1]
port 32 nsew
flabel metal2 9152 0 9180 300 0 FreeSans 240 90 0 0 left_instramp_p_to_gpio5_6[0]
port 33 nsew
flabel metal2 9264 0 9292 300 0 FreeSans 240 90 0 0 left_lp_opamp_n_to_gpio5_5[1]
port 34 nsew
flabel metal2 9376 0 9404 300 0 FreeSans 240 90 0 0 left_lp_opamp_n_to_gpio5_5[0]
port 35 nsew
flabel metal2 9488 0 9516 300 0 FreeSans 240 90 0 0 left_lp_opamp_p_to_gpio5_4[1]
port 36 nsew
flabel metal2 9600 0 9628 300 0 FreeSans 240 90 0 0 left_lp_opamp_p_to_gpio5_4[0]
port 37 nsew
flabel metal2 9712 0 9740 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_n_to_gpio5_3[1]
port 38 nsew
flabel metal2 9824 0 9852 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_n_to_gpio5_3[0]
port 39 nsew
flabel metal2 9936 0 9964 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_p_to_gpio5_2[1]
port 40 nsew
flabel metal2 10048 0 10076 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_p_to_gpio5_2[0]
port 41 nsew
flabel metal2 10160 0 10188 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_n_to_gpio5_1[1]
port 42 nsew
flabel metal2 10272 0 10300 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_n_to_gpio5_1[0]
port 43 nsew
flabel metal2 10384 0 10412 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_p_to_gpio5_0[1]
port 44 nsew
flabel metal2 10496 0 10524 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_p_to_gpio5_0[0]
port 45 nsew
flabel metal2 10608 0 10636 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_gpio4_7[1]
port 46 nsew
flabel metal2 10720 0 10748 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_gpio4_7[0]
port 47 nsew
flabel metal2 10832 0 10860 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_gpio4_6[1]
port 48 nsew
flabel metal2 10944 0 10972 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_gpio4_6[0]
port 49 nsew
flabel metal2 11056 0 11084 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_gpio4_5[1]
port 50 nsew
flabel metal2 11168 0 11196 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_gpio4_5[0]
port 51 nsew
flabel metal2 11280 0 11308 300 0 FreeSans 240 90 0 0 left_instramp_to_gpio4_4[1]
port 52 nsew
flabel metal2 11392 0 11420 300 0 FreeSans 240 90 0 0 left_instramp_to_gpio4_4[0]
port 53 nsew
flabel metal2 11728 0 11756 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_gpio4_3[1]
port 56 nsew
flabel metal2 11840 0 11868 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_gpio4_3[0]
port 57 nsew
flabel metal2 11952 0 11980 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_gpio4_2[1]
port 58 nsew
flabel metal2 12064 0 12092 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_gpio4_2[0]
port 59 nsew
flabel metal2 12176 0 12204 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_gpio4_1[1]
port 60 nsew
flabel metal2 12288 0 12316 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_gpio4_1[0]
port 61 nsew
flabel metal2 12400 0 12428 300 0 FreeSans 240 90 0 0 left_lp_opamp_to_gpio4_0[1]
port 62 nsew
flabel metal2 12512 0 12540 300 0 FreeSans 240 90 0 0 left_lp_opamp_to_gpio4_0[0]
port 63 nsew
flabel metal2 12624 0 12652 300 0 FreeSans 240 90 0 0 left_instramp_to_ulpcomp_p[1]
port 64 nsew
flabel metal2 12736 0 12764 300 0 FreeSans 240 90 0 0 left_instramp_to_ulpcomp_p[0]
port 65 nsew
flabel metal2 12848 0 12876 300 0 FreeSans 240 90 0 0 left_instramp_to_comp_p[1]
port 66 nsew
flabel metal2 12960 0 12988 300 0 FreeSans 240 90 0 0 left_instramp_to_comp_p[0]
port 67 nsew
flabel metal2 13072 0 13100 300 0 FreeSans 240 90 0 0 left_instramp_to_adc0[1]
port 68 nsew
flabel metal2 13184 0 13212 300 0 FreeSans 240 90 0 0 left_instramp_to_adc0[0]
port 69 nsew
flabel metal2 13296 0 13324 300 0 FreeSans 240 90 0 0 left_instramp_to_analog1[1]
port 70 nsew
flabel metal2 13408 0 13436 300 0 FreeSans 240 90 0 0 left_instramp_to_analog1[0]
port 71 nsew
flabel metal2 13520 0 13548 300 0 FreeSans 240 90 0 0 left_instramp_to_amuxbusB[1]
port 72 nsew
flabel metal2 13632 0 13660 300 0 FreeSans 240 90 0 0 left_instramp_to_amuxbusB[0]
port 73 nsew
flabel metal2 13744 0 13772 300 0 FreeSans 240 90 0 0 left_instramp_n_to_analog1
port 74 nsew
flabel metal2 13856 0 13884 300 0 FreeSans 240 90 0 0 left_instramp_n_to_amuxbusB
port 75 nsew
flabel metal2 13968 0 13996 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_ulpcomp_p[1]
port 76 nsew
flabel metal2 14080 0 14108 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_ulpcomp_p[0]
port 77 nsew
flabel metal2 14192 0 14220 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_comp_p[1]
port 78 nsew
flabel metal2 14304 0 14332 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_comp_p[0]
port 79 nsew
flabel metal2 14416 0 14444 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_adc0[1]
port 80 nsew
flabel metal2 14528 0 14556 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_adc0[0]
port 81 nsew
flabel metal2 14640 0 14668 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_ulpcomp_n[1]
port 82 nsew
flabel metal2 14752 0 14780 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_ulpcomp_n[0]
port 83 nsew
flabel metal2 14864 0 14892 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_comp_n[1]
port 84 nsew
flabel metal2 14976 0 15004 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_comp_n[0]
port 85 nsew
flabel metal2 15088 0 15116 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_adc1[1]
port 86 nsew
flabel metal2 15200 0 15228 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_adc1[0]
port 87 nsew
flabel metal2 15312 0 15340 300 0 FreeSans 240 90 0 0 right_instramp_to_ulpcomp_n[1]
port 88 nsew
flabel metal2 15424 0 15452 300 0 FreeSans 240 90 0 0 right_instramp_to_ulpcomp_n[0]
port 89 nsew
flabel metal2 15536 0 15564 300 0 FreeSans 240 90 0 0 right_instramp_to_comp_n[1]
port 90 nsew
flabel metal2 15648 0 15676 300 0 FreeSans 240 90 0 0 right_instramp_to_comp_n[0]
port 91 nsew
flabel metal2 15760 0 15788 300 0 FreeSans 240 90 0 0 right_instramp_to_adc1[1]
port 92 nsew
flabel metal2 15872 0 15900 300 0 FreeSans 240 90 0 0 right_instramp_to_adc1[0]
port 93 nsew
flabel metal2 15984 0 16012 300 0 FreeSans 240 90 0 0 left_instramp_p_to_analog0
port 94 nsew
flabel metal2 16096 0 16124 300 0 FreeSans 240 90 0 0 left_instramp_p_to_amuxbusA
port 95 nsew
flabel metal2 16208 0 16236 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_ulpcomp_p[1]
port 96 nsew
flabel metal2 16320 0 16348 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_ulpcomp_p[0]
port 97 nsew
flabel metal2 16432 0 16460 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_comp_p[1]
port 98 nsew
flabel metal2 16544 0 16572 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_comp_p[0]
port 99 nsew
flabel metal2 16656 0 16684 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_adc0[1]
port 100 nsew
flabel metal2 16768 0 16796 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_adc0[0]
port 101 nsew
flabel metal2 16880 0 16908 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_analog1[1]
port 102 nsew
flabel metal2 16992 0 17020 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_analog1[0]
port 103 nsew
flabel metal2 17104 0 17132 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_amuxbusB[1]
port 104 nsew
flabel metal2 17216 0 17244 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_amuxbusB[0]
port 105 nsew
flabel metal2 17328 0 17356 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_p_to_dac0
port 106 nsew
flabel metal2 17440 0 17468 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_p_to_analog0
port 107 nsew
flabel metal2 17552 0 17580 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_p_to_amuxbusA
port 108 nsew
flabel metal2 17776 0 17804 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_n_to_dac1
port 110 nsew
flabel metal2 17888 0 17916 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_n_to_analog1
port 111 nsew
flabel metal2 18000 0 18028 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_n_to_amuxbusB
port 112 nsew
flabel metal2 18224 0 18252 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_n_to_rheostat_tap
port 114 nsew
flabel metal2 18336 0 18364 300 0 FreeSans 240 90 0 0 left_lp_opamp_to_ulpcomp_n[1]
port 115 nsew
flabel metal2 18448 0 18476 300 0 FreeSans 240 90 0 0 left_lp_opamp_to_ulpcomp_n[0]
port 116 nsew
flabel metal2 18560 0 18588 300 0 FreeSans 240 90 0 0 left_lp_opamp_to_comp_n[1]
port 117 nsew
flabel metal2 18672 0 18700 300 0 FreeSans 240 90 0 0 left_lp_opamp_to_comp_n[0]
port 118 nsew
flabel metal2 18896 0 18924 300 0 FreeSans 240 90 0 0 left_lp_opamp_to_adc1[0]
port 120 nsew
flabel metal2 19008 0 19036 300 0 FreeSans 240 90 0 0 left_lp_opamp_to_analog0[1]
port 121 nsew
flabel metal2 19120 0 19148 300 0 FreeSans 240 90 0 0 left_lp_opamp_to_analog0[0]
port 122 nsew
flabel metal2 19232 0 19260 300 0 FreeSans 240 90 0 0 left_lp_opamp_to_amuxbusA[1]
port 123 nsew
flabel metal2 19344 0 19372 300 0 FreeSans 240 90 0 0 left_lp_opamp_to_amuxbusA[0]
port 124 nsew
flabel metal2 19456 0 19484 300 0 FreeSans 240 90 0 0 left_lp_opamp_p_to_dac0
port 125 nsew
flabel metal2 19568 0 19596 300 0 FreeSans 240 90 0 0 left_lp_opamp_p_to_analog0
port 126 nsew
flabel metal2 19680 0 19708 300 0 FreeSans 240 90 0 0 left_lp_opamp_p_to_amuxbusA
port 127 nsew
flabel metal2 19904 0 19932 300 0 FreeSans 240 90 0 0 left_lp_opamp_n_to_dac1
port 129 nsew
flabel metal2 20016 0 20044 300 0 FreeSans 240 90 0 0 left_lp_opamp_n_to_analog1
port 130 nsew
flabel metal2 20128 0 20156 300 0 FreeSans 240 90 0 0 left_lp_opamp_n_to_amuxbusB
port 131 nsew
flabel metal2 20352 0 20380 300 0 FreeSans 240 90 0 0 left_lp_opamp_n_to_rheostat_tap
port 133 nsew
flabel metal2 527856 0 527884 300 0 FreeSans 240 90 0 0 comp_out
port 244 nsew
flabel metal2 527968 0 527996 300 0 FreeSans 240 90 0 0 ulpcomp_out
port 245 nsew
flabel metal2 528080 0 528108 300 0 FreeSans 240 90 0 0 overvoltage_out
port 246 nsew
flabel metal2 528192 0 528220 300 0 FreeSans 240 90 0 0 comp_ena
port 247 nsew
flabel metal2 528304 0 528332 300 0 FreeSans 240 90 0 0 comp_trim[5]
port 248 nsew
flabel metal2 528416 0 528444 300 0 FreeSans 240 90 0 0 comp_trim[4]
port 249 nsew
flabel metal2 528528 0 528556 300 0 FreeSans 240 90 0 0 comp_trim[3]
port 250 nsew
flabel metal2 528640 0 528668 300 0 FreeSans 240 90 0 0 comp_trim[2]
port 251 nsew
flabel metal2 528752 0 528780 300 0 FreeSans 240 90 0 0 comp_trim[1]
port 252 nsew
flabel metal2 528864 0 528892 300 0 FreeSans 240 90 0 0 comp_trim[0]
port 253 nsew
flabel metal2 528976 0 529004 300 0 FreeSans 240 90 0 0 comp_hyst[1]
port 254 nsew
flabel metal2 529088 0 529116 300 0 FreeSans 240 90 0 0 comp_hyst[0]
port 255 nsew
flabel metal2 529200 0 529228 300 0 FreeSans 240 90 0 0 ulpcomp_ena
port 256 nsew
flabel metal2 529312 0 529340 300 0 FreeSans 240 90 0 0 ulpcomp_clk
port 257 nsew
flabel metal2 529424 0 529452 300 0 FreeSans 240 90 0 0 bandgap_ena
port 258 nsew
flabel metal2 529536 0 529564 300 0 FreeSans 240 90 0 0 bandgap_trim[15]
port 259 nsew
flabel metal2 529648 0 529676 300 0 FreeSans 240 90 0 0 bandgap_trim[14]
port 260 nsew
flabel metal2 529760 0 529788 300 0 FreeSans 240 90 0 0 bandgap_trim[13]
port 261 nsew
flabel metal2 529872 0 529900 300 0 FreeSans 240 90 0 0 bandgap_trim[12]
port 262 nsew
flabel metal2 529984 0 530012 300 0 FreeSans 240 90 0 0 bandgap_trim[11]
port 263 nsew
flabel metal2 530096 0 530124 300 0 FreeSans 240 90 0 0 bandgap_trim[10]
port 264 nsew
flabel metal2 530208 0 530236 300 0 FreeSans 240 90 0 0 bandgap_trim[9]
port 265 nsew
flabel metal2 530320 0 530348 300 0 FreeSans 240 90 0 0 bandgap_trim[8]
port 266 nsew
flabel metal2 530432 0 530460 300 0 FreeSans 240 90 0 0 bandgap_trim[7]
port 267 nsew
flabel metal2 530544 0 530572 300 0 FreeSans 240 90 0 0 bandgap_trim[6]
port 268 nsew
flabel metal2 530656 0 530684 300 0 FreeSans 240 90 0 0 bandgap_trim[5]
port 269 nsew
flabel metal2 530768 0 530796 300 0 FreeSans 240 90 0 0 bandgap_trim[4]
port 270 nsew
flabel metal2 530880 0 530908 300 0 FreeSans 240 90 0 0 bandgap_trim[3]
port 271 nsew
flabel metal2 530992 0 531020 300 0 FreeSans 240 90 0 0 bandgap_trim[2]
port 272 nsew
flabel metal2 531104 0 531132 300 0 FreeSans 240 90 0 0 bandgap_trim[1]
port 273 nsew
flabel metal2 531216 0 531244 300 0 FreeSans 240 90 0 0 bandgap_trim[0]
port 274 nsew
flabel metal2 531328 0 531356 300 0 FreeSans 240 90 0 0 ldo_ena
port 275 nsew
flabel metal2 531440 0 531468 300 0 FreeSans 240 90 0 0 ibias_ena
port 276 nsew
flabel metal2 531552 0 531580 300 0 FreeSans 240 90 0 0 ibias_src_ena[23]
port 277 nsew
flabel metal2 531664 0 531692 300 0 FreeSans 240 90 0 0 ibias_src_ena[22]
port 278 nsew
flabel metal2 531776 0 531804 300 0 FreeSans 240 90 0 0 ibias_src_ena[21]
port 279 nsew
flabel metal2 531888 0 531916 300 0 FreeSans 240 90 0 0 ibias_src_ena[20]
port 280 nsew
flabel metal2 532000 0 532028 300 0 FreeSans 240 90 0 0 ibias_src_ena[19]
port 281 nsew
flabel metal2 532112 0 532140 300 0 FreeSans 240 90 0 0 ibias_src_ena[18]
port 282 nsew
flabel metal2 532224 0 532252 300 0 FreeSans 240 90 0 0 ibias_src_ena[17]
port 283 nsew
flabel metal2 532336 0 532364 300 0 FreeSans 240 90 0 0 ibias_src_ena[16]
port 284 nsew
flabel metal2 532448 0 532476 300 0 FreeSans 240 90 0 0 ibias_src_ena[15]
port 285 nsew
flabel metal2 532560 0 532588 300 0 FreeSans 240 90 0 0 ibias_src_ena[14]
port 286 nsew
flabel metal2 532672 0 532700 300 0 FreeSans 240 90 0 0 ibias_src_ena[13]
port 287 nsew
flabel metal2 532784 0 532812 300 0 FreeSans 240 90 0 0 ibias_src_ena[12]
port 288 nsew
flabel metal2 532896 0 532924 300 0 FreeSans 240 90 0 0 ibias_src_ena[11]
port 289 nsew
flabel metal2 533008 0 533036 300 0 FreeSans 240 90 0 0 ibias_src_ena[10]
port 290 nsew
flabel metal2 533120 0 533148 300 0 FreeSans 240 90 0 0 ibias_src_ena[9]
port 291 nsew
flabel metal2 533232 0 533260 300 0 FreeSans 240 90 0 0 ibias_src_ena[8]
port 292 nsew
flabel metal2 533344 0 533372 300 0 FreeSans 240 90 0 0 ibias_src_ena[7]
port 293 nsew
flabel metal2 533456 0 533484 300 0 FreeSans 240 90 0 0 ibias_src_ena[6]
port 294 nsew
flabel metal2 533568 0 533596 300 0 FreeSans 240 90 0 0 ibias_src_ena[5]
port 295 nsew
flabel metal2 533680 0 533708 300 0 FreeSans 240 90 0 0 ibias_src_ena[4]
port 296 nsew
flabel metal2 533792 0 533820 300 0 FreeSans 240 90 0 0 ibias_src_ena[3]
port 297 nsew
flabel metal2 533904 0 533932 300 0 FreeSans 240 90 0 0 ibias_src_ena[2]
port 298 nsew
flabel metal2 534016 0 534044 300 0 FreeSans 240 90 0 0 ibias_src_ena[1]
port 299 nsew
flabel metal2 534128 0 534156 300 0 FreeSans 240 90 0 0 ibias_src_ena[0]
port 300 nsew
flabel metal2 534240 0 534268 300 0 FreeSans 240 90 0 0 ibias_snk_ena[3]
port 301 nsew
flabel metal2 534352 0 534380 300 0 FreeSans 240 90 0 0 ibias_snk_ena[2]
port 302 nsew
flabel metal2 534464 0 534492 300 0 FreeSans 240 90 0 0 ibias_snk_ena[1]
port 303 nsew
flabel metal2 534576 0 534604 300 0 FreeSans 240 90 0 0 ibias_snk_ena[0]
port 304 nsew
flabel metal2 534688 0 534716 300 0 FreeSans 240 90 0 0 ibias_ref_select
port 305 nsew
flabel metal2 534800 0 534828 300 0 FreeSans 240 90 0 0 overvoltage_ena
port 306 nsew
flabel metal2 534912 0 534940 300 0 FreeSans 240 90 0 0 overvoltage_trim[3]
port 307 nsew
flabel metal2 535024 0 535052 300 0 FreeSans 240 90 0 0 overvoltage_trim[2]
port 308 nsew
flabel metal2 535136 0 535164 300 0 FreeSans 240 90 0 0 overvoltage_trim[1]
port 309 nsew
flabel metal2 535248 0 535276 300 0 FreeSans 240 90 0 0 overvoltage_trim[0]
port 310 nsew
flabel metal2 535360 0 535388 300 0 FreeSans 240 90 0 0 idac_value[11]
port 311 nsew
flabel metal2 535472 0 535500 300 0 FreeSans 240 90 0 0 idac_value[10]
port 312 nsew
flabel metal2 535584 0 535612 300 0 FreeSans 240 90 0 0 idac_value[9]
port 313 nsew
flabel metal2 535696 0 535724 300 0 FreeSans 240 90 0 0 idac_value[8]
port 314 nsew
flabel metal2 535808 0 535836 300 0 FreeSans 240 90 0 0 idac_value[7]
port 315 nsew
flabel metal2 535920 0 535948 300 0 FreeSans 240 90 0 0 idac_value[6]
port 316 nsew
flabel metal2 536032 0 536060 300 0 FreeSans 240 90 0 0 idac_value[5]
port 317 nsew
flabel metal2 536144 0 536172 300 0 FreeSans 240 90 0 0 idac_value[4]
port 318 nsew
flabel metal2 536256 0 536284 300 0 FreeSans 240 90 0 0 idac_value[3]
port 319 nsew
flabel metal2 536368 0 536396 300 0 FreeSans 240 90 0 0 idac_value[2]
port 320 nsew
flabel metal2 536480 0 536508 300 0 FreeSans 240 90 0 0 idac_value[1]
port 321 nsew
flabel metal2 536592 0 536620 300 0 FreeSans 240 90 0 0 idac_value[0]
port 322 nsew
flabel metal2 536704 0 536732 300 0 FreeSans 240 90 0 0 idac_ena
port 323 nsew
flabel metal2 536816 0 536844 300 0 FreeSans 240 90 0 0 right_instramp_ena
port 324 nsew
flabel metal2 536928 0 536956 300 0 FreeSans 240 90 0 0 right_instramp_G1[4]
port 325 nsew
flabel metal2 537040 0 537068 300 0 FreeSans 240 90 0 0 right_instramp_G1[3]
port 326 nsew
flabel metal2 537152 0 537180 300 0 FreeSans 240 90 0 0 right_instramp_G1[2]
port 327 nsew
flabel metal2 537264 0 537292 300 0 FreeSans 240 90 0 0 right_instramp_G1[1]
port 328 nsew
flabel metal2 537376 0 537404 300 0 FreeSans 240 90 0 0 right_instramp_G1[0]
port 329 nsew
flabel metal2 537488 0 537516 300 0 FreeSans 240 90 0 0 right_instramp_G2[4]
port 330 nsew
flabel metal2 537600 0 537628 300 0 FreeSans 240 90 0 0 right_instramp_G2[3]
port 331 nsew
flabel metal2 537712 0 537740 300 0 FreeSans 240 90 0 0 right_instramp_G2[2]
port 332 nsew
flabel metal2 537824 0 537852 300 0 FreeSans 240 90 0 0 right_instramp_G2[1]
port 333 nsew
flabel metal2 537936 0 537964 300 0 FreeSans 240 90 0 0 right_instramp_G2[0]
port 334 nsew
flabel metal2 538048 0 538076 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_ena
port 335 nsew
flabel metal2 538160 0 538188 300 0 FreeSans 240 90 0 0 right_lp_opamp_ena
port 336 nsew
flabel metal2 538272 0 538300 300 0 FreeSans 240 90 0 0 right_rheostat1_b[7]
port 337 nsew
flabel metal2 538384 0 538412 300 0 FreeSans 240 90 0 0 right_rheostat1_b[6]
port 338 nsew
flabel metal2 538496 0 538524 300 0 FreeSans 240 90 0 0 right_rheostat1_b[5]
port 339 nsew
flabel metal2 538608 0 538636 300 0 FreeSans 240 90 0 0 right_rheostat1_b[4]
port 340 nsew
flabel metal2 538720 0 538748 300 0 FreeSans 240 90 0 0 right_rheostat1_b[3]
port 341 nsew
flabel metal2 538832 0 538860 300 0 FreeSans 240 90 0 0 right_rheostat1_b[2]
port 342 nsew
flabel metal2 538944 0 538972 300 0 FreeSans 240 90 0 0 right_rheostat1_b[1]
port 343 nsew
flabel metal2 539056 0 539084 300 0 FreeSans 240 90 0 0 right_rheostat1_b[0]
port 344 nsew
flabel metal2 539168 0 539196 300 0 FreeSans 240 90 0 0 right_rheostat2_b[7]
port 345 nsew
flabel metal2 539280 0 539308 300 0 FreeSans 240 90 0 0 right_rheostat2_b[6]
port 346 nsew
flabel metal2 539392 0 539420 300 0 FreeSans 240 90 0 0 right_rheostat2_b[5]
port 347 nsew
flabel metal2 539504 0 539532 300 0 FreeSans 240 90 0 0 right_rheostat2_b[4]
port 348 nsew
flabel metal2 539616 0 539644 300 0 FreeSans 240 90 0 0 right_rheostat2_b[3]
port 349 nsew
flabel metal2 539728 0 539756 300 0 FreeSans 240 90 0 0 right_rheostat2_b[2]
port 350 nsew
flabel metal2 539840 0 539868 300 0 FreeSans 240 90 0 0 right_rheostat2_b[1]
port 351 nsew
flabel metal2 539952 0 539980 300 0 FreeSans 240 90 0 0 right_rheostat2_b[0]
port 352 nsew
flabel metal2 540064 0 540092 300 0 FreeSans 240 90 0 0 por
port 353 nsew
flabel metal2 540176 0 540204 300 0 FreeSans 240 90 0 0 porb
port 354 nsew
flabel metal2 540400 0 540428 300 0 FreeSans 240 90 0 0 user_to_comp_n[1]
port 356 nsew
flabel metal2 540512 0 540540 300 0 FreeSans 240 90 0 0 user_to_comp_n[0]
port 357 nsew
flabel metal2 540624 0 540652 300 0 FreeSans 240 90 0 0 user_to_comp_p[1]
port 358 nsew
flabel metal2 540736 0 540764 300 0 FreeSans 240 90 0 0 user_to_comp_p[0]
port 359 nsew
flabel metal2 540848 0 540876 300 0 FreeSans 240 90 0 0 user_to_ulpcomp_n[1]
port 360 nsew
flabel metal2 540960 0 540988 300 0 FreeSans 240 90 0 0 user_to_ulpcomp_n[0]
port 361 nsew
flabel metal2 541072 0 541100 300 0 FreeSans 240 90 0 0 user_to_ulpcomp_p[1]
port 362 nsew
flabel metal2 541184 0 541212 300 0 FreeSans 240 90 0 0 user_to_ulpcomp_p[0]
port 363 nsew
flabel metal2 541296 0 541324 300 0 FreeSans 240 90 0 0 user_to_adc0[1]
port 364 nsew
flabel metal2 541408 0 541436 300 0 FreeSans 240 90 0 0 user_to_adc0[0]
port 365 nsew
flabel metal2 541520 0 541548 300 0 FreeSans 240 90 0 0 user_to_adc1[1]
port 366 nsew
flabel metal2 541632 0 541660 300 0 FreeSans 240 90 0 0 user_to_adc1[0]
port 367 nsew
flabel metal2 541744 0 541772 300 0 FreeSans 240 90 0 0 dac0_to_user
port 368 nsew
flabel metal2 541856 0 541884 300 0 FreeSans 240 90 0 0 dac1_to_user
port 369 nsew
flabel metal2 541968 0 541996 300 0 FreeSans 240 90 0 0 tempsense_to_user
port 370 nsew
flabel metal2 542080 0 542108 300 0 FreeSans 240 90 0 0 right_vref_to_user
port 371 nsew
flabel metal2 542192 0 542220 300 0 FreeSans 240 90 0 0 left_vref_to_user
port 372 nsew
flabel metal2 542304 0 542332 300 0 FreeSans 240 90 0 0 vinref_to_user
port 373 nsew
flabel metal2 542416 0 542444 300 0 FreeSans 240 90 0 0 voutref_to_user
port 374 nsew
flabel metal2 542528 0 542556 300 0 FreeSans 240 90 0 0 vbgtc_to_user
port 375 nsew
flabel metal2 542640 0 542668 300 0 FreeSans 240 90 0 0 vbgsc_to_user
port 376 nsew
flabel metal2 542752 0 542780 300 0 FreeSans 240 90 0 0 sio0_connect[1]
port 377 nsew
flabel metal2 542864 0 542892 300 0 FreeSans 240 90 0 0 sio0_connect[0]
port 378 nsew
flabel metal2 542976 0 543004 300 0 FreeSans 240 90 0 0 sio1_connect[1]
port 379 nsew
flabel metal2 543088 0 543116 300 0 FreeSans 240 90 0 0 sio1_connect[0]
port 380 nsew
flabel metal2 543200 0 543228 300 0 FreeSans 240 90 0 0 comp_p_to_dac0
port 381 nsew
flabel metal2 543312 0 543340 300 0 FreeSans 240 90 0 0 comp_p_to_analog1
port 382 nsew
flabel metal2 543424 0 543452 300 0 FreeSans 240 90 0 0 comp_p_to_sio0
port 383 nsew
flabel metal2 543536 0 543564 300 0 FreeSans 240 90 0 0 comp_p_to_vbgtc
port 384 nsew
flabel metal2 543648 0 543676 300 0 FreeSans 240 90 0 0 comp_p_to_tempsense
port 385 nsew
flabel metal2 543760 0 543788 300 0 FreeSans 240 90 0 0 comp_p_to_left_vref
port 386 nsew
flabel metal2 543872 0 543900 300 0 FreeSans 240 90 0 0 comp_p_to_voutref
port 387 nsew
flabel metal2 543984 0 544012 300 0 FreeSans 240 90 0 0 comp_n_to_dac1
port 388 nsew
flabel metal2 544096 0 544124 300 0 FreeSans 240 90 0 0 comp_n_to_analog0
port 389 nsew
flabel metal2 544208 0 544236 300 0 FreeSans 240 90 0 0 comp_n_to_sio1
port 390 nsew
flabel metal2 544320 0 544348 300 0 FreeSans 240 90 0 0 comp_n_to_vbgsc
port 391 nsew
flabel metal2 544432 0 544460 300 0 FreeSans 240 90 0 0 comp_n_to_right_vref
port 392 nsew
flabel metal2 544544 0 544572 300 0 FreeSans 240 90 0 0 comp_n_to_vinref
port 393 nsew
flabel metal2 544656 0 544684 300 0 FreeSans 240 90 0 0 ulpcomp_p_to_dac0
port 394 nsew
flabel metal2 544768 0 544796 300 0 FreeSans 240 90 0 0 ulpcomp_p_to_analog1
port 395 nsew
flabel metal2 544880 0 544908 300 0 FreeSans 240 90 0 0 ulpcomp_p_to_sio0
port 396 nsew
flabel metal2 544992 0 545020 300 0 FreeSans 240 90 0 0 ulpcomp_p_to_vbgtc
port 397 nsew
flabel metal2 545104 0 545132 300 0 FreeSans 240 90 0 0 ulpcomp_p_to_tempsense
port 398 nsew
flabel metal2 545216 0 545244 300 0 FreeSans 240 90 0 0 ulpcomp_p_to_left_vref
port 399 nsew
flabel metal2 545328 0 545356 300 0 FreeSans 240 90 0 0 ulpcomp_p_to_voutref
port 400 nsew
flabel metal2 545440 0 545468 300 0 FreeSans 240 90 0 0 ulpcomp_n_to_dac1
port 401 nsew
flabel metal2 545552 0 545580 300 0 FreeSans 240 90 0 0 ulpcomp_n_to_analog0
port 402 nsew
flabel metal2 545664 0 545692 300 0 FreeSans 240 90 0 0 ulpcomp_n_to_sio1
port 403 nsew
flabel metal2 545776 0 545804 300 0 FreeSans 240 90 0 0 ulpcomp_n_to_vbgsc
port 404 nsew
flabel metal2 545888 0 545916 300 0 FreeSans 240 90 0 0 ulpcomp_n_to_right_vref
port 405 nsew
flabel metal2 546000 0 546028 300 0 FreeSans 240 90 0 0 ulpcomp_n_to_vinref
port 406 nsew
flabel metal2 546112 0 546140 300 0 FreeSans 240 90 0 0 left_instramp_n_to_sio1
port 407 nsew
flabel metal2 546224 0 546252 300 0 FreeSans 240 90 0 0 left_instramp_n_to_right_vref
port 408 nsew
flabel metal2 546336 0 546364 300 0 FreeSans 240 90 0 0 left_instramp_n_to_vinref
port 409 nsew
flabel metal2 546448 0 546476 300 0 FreeSans 240 90 0 0 left_instramp_p_to_sio0
port 410 nsew
flabel metal2 546560 0 546588 300 0 FreeSans 240 90 0 0 left_instramp_p_to_tempsense
port 411 nsew
flabel metal2 546672 0 546700 300 0 FreeSans 240 90 0 0 left_instramp_p_to_left_vref
port 412 nsew
flabel metal2 546784 0 546812 300 0 FreeSans 240 90 0 0 left_instramp_p_to_voutref
port 413 nsew
flabel metal2 546896 0 546924 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_p_to_sio0
port 414 nsew
flabel metal2 547008 0 547036 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_p_to_tempsense
port 415 nsew
flabel metal2 547120 0 547148 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_p_to_left_vref
port 416 nsew
flabel metal2 547232 0 547260 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_p_to_voutref
port 417 nsew
flabel metal2 547344 0 547372 300 0 FreeSans 240 90 0 0 left_lp_opamp_p_to_sio0
port 418 nsew
flabel metal2 547456 0 547484 300 0 FreeSans 240 90 0 0 left_lp_opamp_p_to_left_vref
port 419 nsew
flabel metal2 547568 0 547596 300 0 FreeSans 240 90 0 0 left_lp_opamp_p_to_voutref
port 420 nsew
flabel metal2 547680 0 547708 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_n_to_sio1
port 421 nsew
flabel metal2 547792 0 547820 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_n_to_vbgtc
port 422 nsew
flabel metal2 547904 0 547932 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_n_to_right_vref
port 423 nsew
flabel metal2 548016 0 548044 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_n_to_vinref
port 424 nsew
flabel metal2 548128 0 548156 300 0 FreeSans 240 90 0 0 left_lp_opamp_n_to_sio1
port 425 nsew
flabel metal2 548240 0 548268 300 0 FreeSans 240 90 0 0 left_lp_opamp_n_to_vbgsc
port 426 nsew
flabel metal2 548352 0 548380 300 0 FreeSans 240 90 0 0 left_lp_opamp_n_to_right_vref
port 427 nsew
flabel metal2 548464 0 548492 300 0 FreeSans 240 90 0 0 left_lp_opamp_n_to_vinref
port 428 nsew
flabel metal2 548576 0 548604 300 0 FreeSans 240 90 0 0 adc0_to_vbgtc
port 429 nsew
flabel metal2 548688 0 548716 300 0 FreeSans 240 90 0 0 adc0_to_tempsense
port 430 nsew
flabel metal2 548800 0 548828 300 0 FreeSans 240 90 0 0 adc0_to_left_vref
port 431 nsew
flabel metal2 548912 0 548940 300 0 FreeSans 240 90 0 0 adc0_to_voutref
port 432 nsew
flabel metal2 549024 0 549052 300 0 FreeSans 240 90 0 0 adc1_to_vbgsc
port 433 nsew
flabel metal2 549136 0 549164 300 0 FreeSans 240 90 0 0 adc1_to_right_vref
port 434 nsew
flabel metal2 549248 0 549276 300 0 FreeSans 240 90 0 0 adc1_to_vinref
port 435 nsew
flabel metal2 549360 0 549388 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_analog1[1]
port 436 nsew
flabel metal2 549472 0 549500 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_analog1[0]
port 437 nsew
flabel metal2 549584 0 549612 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_amuxbusB[1]
port 438 nsew
flabel metal2 549696 0 549724 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_amuxbusB[0]
port 439 nsew
flabel metal2 549808 0 549836 300 0 FreeSans 240 90 0 0 right_lp_opamp_p_to_dac0
port 440 nsew
flabel metal2 549920 0 549948 300 0 FreeSans 240 90 0 0 right_lp_opamp_p_to_analog0
port 441 nsew
flabel metal2 550032 0 550060 300 0 FreeSans 240 90 0 0 right_lp_opamp_p_to_amuxbusA
port 442 nsew
flabel metal2 550256 0 550284 300 0 FreeSans 240 90 0 0 right_lp_opamp_p_to_sio0
port 444 nsew
flabel metal2 550368 0 550396 300 0 FreeSans 240 90 0 0 right_lp_opamp_p_to_tempsense
port 445 nsew
flabel metal2 550480 0 550508 300 0 FreeSans 240 90 0 0 right_lp_opamp_p_to_left_vref
port 446 nsew
flabel metal2 550592 0 550620 300 0 FreeSans 240 90 0 0 right_lp_opamp_p_to_voutref
port 447 nsew
flabel metal2 550704 0 550732 300 0 FreeSans 240 90 0 0 right_lp_opamp_n_to_dac1
port 448 nsew
flabel metal2 550816 0 550844 300 0 FreeSans 240 90 0 0 right_lp_opamp_n_to_analog1
port 449 nsew
flabel metal2 550928 0 550956 300 0 FreeSans 240 90 0 0 right_lp_opamp_n_to_amuxbusB
port 450 nsew
flabel metal2 551152 0 551180 300 0 FreeSans 240 90 0 0 right_lp_opamp_n_to_rheostat_tap
port 452 nsew
flabel metal2 551264 0 551292 300 0 FreeSans 240 90 0 0 right_lp_opamp_n_to_sio1
port 453 nsew
flabel metal2 551376 0 551404 300 0 FreeSans 240 90 0 0 right_lp_opamp_n_to_vbgtc
port 454 nsew
flabel metal2 551488 0 551516 300 0 FreeSans 240 90 0 0 right_lp_opamp_n_to_right_vref
port 455 nsew
flabel metal2 551600 0 551628 300 0 FreeSans 240 90 0 0 right_lp_opamp_n_to_vinref
port 456 nsew
flabel metal2 551712 0 551740 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_analog0[1]
port 457 nsew
flabel metal2 551824 0 551852 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_analog0[0]
port 458 nsew
flabel metal2 551936 0 551964 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_amuxbusA[1]
port 459 nsew
flabel metal2 552048 0 552076 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_amuxbusA[0]
port 460 nsew
flabel metal2 552160 0 552188 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_p_to_dac0
port 461 nsew
flabel metal2 552272 0 552300 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_p_to_analog0
port 462 nsew
flabel metal2 552384 0 552412 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_p_to_amuxbusA
port 463 nsew
flabel metal2 552608 0 552636 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_p_to_sio0
port 465 nsew
flabel metal2 552720 0 552748 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_p_to_left_vref
port 466 nsew
flabel metal2 552832 0 552860 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_p_to_voutref
port 467 nsew
flabel metal2 552944 0 552972 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_n_to_dac1
port 468 nsew
flabel metal2 553056 0 553084 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_n_to_analog1
port 469 nsew
flabel metal2 553168 0 553196 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_n_to_amuxbusB
port 470 nsew
flabel metal2 553392 0 553420 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_n_to_rheostat_tap
port 472 nsew
flabel metal2 553504 0 553532 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_n_to_sio1
port 473 nsew
flabel metal2 553616 0 553644 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_n_to_vbgsc
port 474 nsew
flabel metal2 553728 0 553756 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_n_to_right_vref
port 475 nsew
flabel metal2 553840 0 553868 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_n_to_vinref
port 476 nsew
flabel metal2 553952 0 553980 300 0 FreeSans 240 90 0 0 right_instramp_to_analog0[1]
port 477 nsew
flabel metal2 554064 0 554092 300 0 FreeSans 240 90 0 0 right_instramp_to_analog0[0]
port 478 nsew
flabel metal2 554176 0 554204 300 0 FreeSans 240 90 0 0 right_instramp_to_amuxbusA[1]
port 479 nsew
flabel metal2 554288 0 554316 300 0 FreeSans 240 90 0 0 right_instramp_to_amuxbusA[0]
port 480 nsew
flabel metal2 554400 0 554428 300 0 FreeSans 240 90 0 0 right_instramp_n_to_analog1
port 481 nsew
flabel metal2 554512 0 554540 300 0 FreeSans 240 90 0 0 right_instramp_n_to_amuxbusB
port 482 nsew
flabel metal2 554624 0 554652 300 0 FreeSans 240 90 0 0 right_instramp_n_to_sio1
port 483 nsew
flabel metal2 554736 0 554764 300 0 FreeSans 240 90 0 0 right_instramp_n_to_right_vref
port 484 nsew
flabel metal2 554848 0 554876 300 0 FreeSans 240 90 0 0 right_instramp_n_to_vinref
port 485 nsew
flabel metal2 554960 0 554988 300 0 FreeSans 240 90 0 0 right_instramp_p_to_analog0
port 486 nsew
flabel metal2 555072 0 555100 300 0 FreeSans 240 90 0 0 right_instramp_p_to_amuxbusA
port 487 nsew
flabel metal2 555184 0 555212 300 0 FreeSans 240 90 0 0 right_instramp_p_to_tempsense
port 488 nsew
flabel metal2 555296 0 555324 300 0 FreeSans 240 90 0 0 right_instramp_p_to_left_vref
port 489 nsew
flabel metal2 555408 0 555436 300 0 FreeSans 240 90 0 0 right_instramp_p_to_voutref
port 490 nsew
flabel metal2 555520 0 555548 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_gpio3_7[1]
port 491 nsew
flabel metal2 555632 0 555660 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_gpio3_7[0]
port 492 nsew
flabel metal2 555744 0 555772 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_gpio3_6[1]
port 493 nsew
flabel metal2 555856 0 555884 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_gpio3_6[0]
port 494 nsew
flabel metal2 555968 0 555996 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_gpio3_5[1]
port 495 nsew
flabel metal2 556080 0 556108 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_gpio3_5[0]
port 496 nsew
flabel metal2 556192 0 556220 300 0 FreeSans 240 90 0 0 left_lp_opamp_to_gpio3_4[1]
port 497 nsew
flabel metal2 556304 0 556332 300 0 FreeSans 240 90 0 0 left_lp_opamp_to_gpio3_4[0]
port 498 nsew
flabel metal2 556416 0 556444 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_gpio3_3[1]
port 499 nsew
flabel metal2 556528 0 556556 300 0 FreeSans 240 90 0 0 right_lp_opamp_to_gpio3_3[0]
port 500 nsew
flabel metal2 556640 0 556668 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_gpio3_2[1]
port 501 nsew
flabel metal2 556752 0 556780 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_to_gpio3_2[0]
port 502 nsew
flabel metal2 556864 0 556892 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_gpio3_1[1]
port 503 nsew
flabel metal2 556976 0 557004 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_to_gpio3_1[0]
port 504 nsew
flabel metal2 557088 0 557116 300 0 FreeSans 240 90 0 0 right_instramp_to_gpio3_0[1]
port 505 nsew
flabel metal2 557200 0 557228 300 0 FreeSans 240 90 0 0 right_instramp_to_gpio3_0[0]
port 506 nsew
flabel metal2 557536 0 557564 300 0 FreeSans 240 90 0 0 right_instramp_p_to_gpio2_7[1]
port 509 nsew
flabel metal2 557648 0 557676 300 0 FreeSans 240 90 0 0 right_instramp_p_to_gpio2_7[0]
port 510 nsew
flabel metal2 557760 0 557788 300 0 FreeSans 240 90 0 0 right_instramp_n_to_gpio2_6[1]
port 511 nsew
flabel metal2 557872 0 557900 300 0 FreeSans 240 90 0 0 right_instramp_n_to_gpio2_6[0]
port 512 nsew
flabel metal2 557984 0 558012 300 0 FreeSans 240 90 0 0 right_lp_opamp_p_to_gpio2_5[1]
port 513 nsew
flabel metal2 558096 0 558124 300 0 FreeSans 240 90 0 0 right_lp_opamp_p_to_gpio2_5[0]
port 514 nsew
flabel metal2 558208 0 558236 300 0 FreeSans 240 90 0 0 right_lp_opamp_n_to_gpio2_4[1]
port 515 nsew
flabel metal2 558320 0 558348 300 0 FreeSans 240 90 0 0 right_lp_opamp_n_to_gpio2_4[0]
port 516 nsew
flabel metal2 558432 0 558460 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_p_to_gpio2_3[1]
port 517 nsew
flabel metal2 558544 0 558572 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_p_to_gpio2_3[0]
port 518 nsew
flabel metal2 558656 0 558684 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_n_to_gpio2_2[1]
port 519 nsew
flabel metal2 558768 0 558796 300 0 FreeSans 240 90 0 0 right_hgbw_opamp_n_to_gpio2_2[0]
port 520 nsew
flabel metal2 558880 0 558908 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_p_to_gpio2_1[1]
port 521 nsew
flabel metal2 558992 0 559020 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_p_to_gpio2_1[0]
port 522 nsew
flabel metal2 559104 0 559132 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_n_to_gpio2_0[1]
port 523 nsew
flabel metal2 559216 0 559244 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_n_to_gpio2_0[0]
port 524 nsew
flabel metal2 559328 0 559356 300 0 FreeSans 240 90 0 0 ulpcomp_p_to_gpio1_7[1]
port 525 nsew
flabel metal2 559440 0 559468 300 0 FreeSans 240 90 0 0 ulpcomp_p_to_gpio1_7[0]
port 526 nsew
flabel metal2 559552 0 559580 300 0 FreeSans 240 90 0 0 ulpcomp_n_to_gpio1_6[1]
port 527 nsew
flabel metal2 559664 0 559692 300 0 FreeSans 240 90 0 0 ulpcomp_n_to_gpio1_6[0]
port 528 nsew
flabel metal2 559776 0 559804 300 0 FreeSans 240 90 0 0 comp_p_to_gpio1_5[1]
port 529 nsew
flabel metal2 559888 0 559916 300 0 FreeSans 240 90 0 0 comp_p_to_gpio1_5[0]
port 530 nsew
flabel metal2 560000 0 560028 300 0 FreeSans 240 90 0 0 comp_n_to_gpio1_4[1]
port 531 nsew
flabel metal2 560112 0 560140 300 0 FreeSans 240 90 0 0 comp_n_to_gpio1_4[0]
port 532 nsew
flabel metal2 560224 0 560252 300 0 FreeSans 240 90 0 0 adc0_to_gpio1_3[1]
port 533 nsew
flabel metal2 560336 0 560364 300 0 FreeSans 240 90 0 0 adc0_to_gpio1_3[0]
port 534 nsew
flabel metal2 560448 0 560476 300 0 FreeSans 240 90 0 0 idac_to_gpio1_3[1]
port 535 nsew
flabel metal2 560560 0 560588 300 0 FreeSans 240 90 0 0 idac_to_gpio1_3[0]
port 536 nsew
flabel metal2 560672 0 560700 300 0 FreeSans 240 90 0 0 ibias_test_to_gpio1_2[1]
port 537 nsew
flabel metal2 560784 0 560812 300 0 FreeSans 240 90 0 0 ibias_test_to_gpio1_2[0]
port 538 nsew
flabel metal2 560896 0 560924 300 0 FreeSans 240 90 0 0 idac_to_gpio1_2[1]
port 539 nsew
flabel metal2 561008 0 561036 300 0 FreeSans 240 90 0 0 idac_to_gpio1_2[0]
port 540 nsew
flabel metal2 561120 0 561148 300 0 FreeSans 240 90 0 0 adc1_to_gpio1_2[1]
port 541 nsew
flabel metal2 561232 0 561260 300 0 FreeSans 240 90 0 0 adc1_to_gpio1_2[0]
port 542 nsew
flabel metal2 561344 0 561372 300 0 FreeSans 240 90 0 0 dac_refh_to_gpio1_1[1]
port 543 nsew
flabel metal2 561456 0 561484 300 0 FreeSans 240 90 0 0 dac_refh_to_gpio1_1[0]
port 544 nsew
flabel metal2 561568 0 561596 300 0 FreeSans 240 90 0 0 vbg_test_to_gpio1_1[1]
port 545 nsew
flabel metal2 561680 0 561708 300 0 FreeSans 240 90 0 0 vbg_test_to_gpio1_1[0]
port 546 nsew
flabel metal5 0 29220 300 29540 0 FreeSans 480 0 0 0 gpio5_3
port 569 nsew
flabel metal5 0 50220 300 50540 0 FreeSans 480 0 0 0 gpio5_2
port 570 nsew
flabel metal5 0 71220 300 71540 0 FreeSans 480 0 0 0 gpio5_1
port 571 nsew
flabel metal5 0 92220 300 92540 0 FreeSans 480 0 0 0 gpio5_0
port 572 nsew
flabel metal5 574300 13200 574600 13520 0 FreeSans 800 0 0 0 gpio2_4
port 593 nsew
flabel metal5 574300 34200 574600 34520 0 FreeSans 800 0 0 0 gpio2_5
port 594 nsew
flabel metal5 574300 55200 574600 55520 0 FreeSans 800 0 0 0 gpio2_6
port 595 nsew
flabel metal5 574300 76200 574600 76520 0 FreeSans 800 0 0 0 gpio2_7
port 596 nsew
flabel metal5 -6 4557 514 9557 0 FreeSans 4000 90 0 0 vdda2
port 597 nsew
flabel metal5 -6 11557 514 16557 0 FreeSans 4000 90 0 0 vssa2
port 598 nsew
flabel metal4 297812 114900 298012 115200 0 FreeSans 480 90 0 0 amuxbus_a_n
port 584 nsew
flabel metal4 297012 114900 297212 115200 0 FreeSans 480 90 0 0 amuxbus_b_n
port 583 nsew
flabel metal4 288812 114900 289012 115200 0 FreeSans 480 90 0 0 analog0
port 582 nsew
flabel metal4 265812 114900 266012 115200 0 FreeSans 480 90 0 0 analog1
port 581 nsew
flabel metal4 222812 114900 223012 115200 0 FreeSans 480 90 0 0 gpio4_0
port 580 nsew
flabel metal4 198812 114900 199012 115200 0 FreeSans 480 90 0 0 gpio4_1
port 579 nsew
flabel metal4 174812 114900 175012 115200 0 FreeSans 480 90 0 0 gpio4_2
port 578 nsew
flabel metal4 150812 114900 151012 115200 0 FreeSans 480 90 0 0 gpio4_3
port 577 nsew
flabel metal4 56812 114900 57012 115200 0 FreeSans 480 90 0 0 gpio4_5
port 575 nsew
flabel metal4 32812 114900 33012 115200 0 FreeSans 480 90 0 0 gpio4_6
port 574 nsew
flabel metal4 8812 114900 9012 115200 0 FreeSans 480 90 0 0 gpio4_7
port 573 nsew
flabel metal4 569700 114900 569900 115200 0 FreeSans 480 90 0 0 gpio3_0
port 592 nsew
flabel metal4 551812 114900 552012 115200 0 FreeSans 480 90 0 0 gpio3_1
port 591 nsew
flabel metal4 527812 114900 528012 115200 0 FreeSans 480 90 0 0 gpio3_2
port 590 nsew
flabel metal4 433812 114900 434012 115200 0 FreeSans 480 90 0 0 gpio3_4
port 588 nsew
flabel metal4 409812 114900 410012 115200 0 FreeSans 480 90 0 0 gpio3_5
port 587 nsew
flabel metal4 385812 114900 386012 115200 0 FreeSans 480 90 0 0 gpio3_6
port 586 nsew
flabel metal4 361812 114900 362012 115200 0 FreeSans 480 90 0 0 gpio3_7
port 585 nsew
flabel metal4 346256 0 346384 300 0 FreeSans 240 90 0 0 user_voutref
port 213 nsew
flabel metal4 346768 0 346896 300 0 FreeSans 240 90 0 0 user_vinref
port 214 nsew
flabel metal4 347280 0 347408 300 0 FreeSans 240 90 0 0 user_left_vref
port 215 nsew
flabel metal4 347792 0 347920 300 0 FreeSans 240 90 0 0 user_right_vref
port 216 nsew
flabel metal4 348304 0 348432 300 0 FreeSans 240 90 0 0 user_tempsense
port 217 nsew
flabel metal4 348816 0 348944 300 0 FreeSans 240 90 0 0 user_dac0
port 218 nsew
flabel metal4 349328 0 349456 300 0 FreeSans 240 90 0 0 user_dac1
port 219 nsew
flabel metal4 349840 0 349968 300 0 FreeSans 240 90 0 0 user_vbgtc
port 220 nsew
flabel metal4 350352 0 350480 300 0 FreeSans 240 90 0 0 user_vbgsc
port 221 nsew
flabel metal4 563952 0 564080 300 0 FreeSans 240 90 0 0 voutref
port 553 nsew
flabel metal4 563440 0 563568 300 0 FreeSans 240 90 0 0 vinref
port 554 nsew
flabel metal4 564464 0 564592 300 0 FreeSans 240 90 0 0 vbg
port 555 nsew
flabel metal4 564976 0 565104 300 0 FreeSans 240 90 0 0 sio0
port 551 nsew
flabel metal4 565488 0 565616 300 0 FreeSans 240 90 0 0 sio1
port 552 nsew
flabel metal4 562928 0 563056 300 0 FreeSans 240 90 0 0 ibias_lsxo
port 549 nsew
flabel metal4 562416 0 562544 300 0 FreeSans 240 90 0 0 ibias_hsxo
port 550 nsew
flabel metal4 351888 0 352016 300 0 FreeSans 240 90 0 0 user_adc0
port 222 nsew
flabel metal4 352400 0 352528 300 0 FreeSans 240 90 0 0 user_adc1
port 223 nsew
flabel metal4 352912 0 353040 300 0 FreeSans 240 90 0 0 user_comp_n
port 224 nsew
flabel metal4 353424 0 353552 300 0 FreeSans 240 90 0 0 user_comp_p
port 225 nsew
flabel metal4 353936 0 354064 300 0 FreeSans 240 90 0 0 user_ulpcomp_n
port 226 nsew
flabel metal4 354448 0 354576 300 0 FreeSans 240 90 0 0 user_ulpcomp_p
port 227 nsew
flabel metal4 354960 0 355088 300 0 FreeSans 240 90 0 0 user_gpio4_7_analog
port 228 nsew
flabel metal4 355472 0 355600 300 0 FreeSans 240 90 0 0 user_gpio4_6_analog
port 229 nsew
flabel metal4 355984 0 356112 300 0 FreeSans 240 90 0 0 user_gpio4_5_analog
port 230 nsew
flabel metal4 356496 0 356624 300 0 FreeSans 240 90 0 0 user_gpio4_4_analog
port 231 nsew
flabel metal4 357008 0 357136 300 0 FreeSans 240 90 0 0 user_gpio4_3_analog
port 232 nsew
flabel metal4 357520 0 357648 300 0 FreeSans 240 90 0 0 user_gpio4_2_analog
port 233 nsew
flabel metal4 358032 0 358160 300 0 FreeSans 240 90 0 0 user_gpio4_1_analog
port 234 nsew
flabel metal4 358544 0 358672 300 0 FreeSans 240 90 0 0 user_gpio4_0_analog
port 235 nsew
flabel metal4 359056 0 359184 300 0 FreeSans 240 90 0 0 user_gpio3_7_analog
port 236 nsew
flabel metal4 359568 0 359696 300 0 FreeSans 240 90 0 0 user_gpio3_6_analog
port 237 nsew
flabel metal4 360080 0 360208 300 0 FreeSans 240 90 0 0 user_gpio3_5_analog
port 238 nsew
flabel metal4 360592 0 360720 300 0 FreeSans 240 90 0 0 user_gpio3_4_analog
port 239 nsew
flabel metal4 361104 0 361232 300 0 FreeSans 240 90 0 0 user_gpio3_3_analog
port 240 nsew
flabel metal4 361616 0 361744 300 0 FreeSans 240 90 0 0 user_gpio3_2_analog
port 241 nsew
flabel metal4 362128 0 362256 300 0 FreeSans 240 90 0 0 user_gpio3_1_analog
port 242 nsew
flabel metal4 362640 0 362768 300 0 FreeSans 240 90 0 0 user_gpio3_0_analog
port 243 nsew
flabel metal4 350864 0 350992 300 0 FreeSans 240 90 0 0 user_ibias50
port 605 nsew
flabel metal4 351376 0 351504 300 0 FreeSans 240 90 0 0 user_ibias100
port 606 nsew
flabel comment s 284054 112372 284054 112372 0 FreeSans 960 90 0 0 analog0
flabel comment s 283244 112340 283244 112340 0 FreeSans 960 90 0 0 analog1
flabel metal5 574084 25557 574604 30557 0 FreeSans 4000 270 0 0 vdda1
port 604 nsew
flabel metal5 574084 18557 574604 23557 0 FreeSans 4000 270 0 0 vssa1
port 603 nsew
flabel metal4 120452 114792 125328 115192 0 FreeSans 3200 0 0 0 vccd2
port 599 nsew
flabel metal4 115352 114792 120228 115192 0 FreeSans 3200 0 0 0 vssd2
port 600 nsew
flabel metal4 303318 114800 308118 115200 0 FreeSans 1600 0 0 0 vdda0
port 607 nsew
flabel metal4 313018 114800 317818 115200 0 FreeSans 1600 0 0 0 vdda0
port 607 nsew
flabel metal4 445288 114800 450164 115200 0 FreeSans 3200 0 0 0 vccd1
port 602 nsew
flabel metal4 450478 114800 455172 115200 0 FreeSans 3200 0 0 0 vssd1
port 601 nsew
flabel metal4 244018 114800 248818 115200 0 FreeSans 1600 0 0 0 vssa0
port 608 nsew
flabel metal4 234318 114800 239118 115200 0 FreeSans 1600 0 0 0 vssa0
port 608 nsew
flabel metal2 527744 0 527772 300 0 FreeSans 240 90 0 0 bandgap_sel
port 612 nsew
flabel metal2 527632 0 527660 300 0 FreeSans 240 90 0 0 ldo_ref_sel
port 613 nsew
flabel metal2 527520 0 527548 300 0 FreeSans 240 90 0 0 tempsense_sel
port 614 nsew
flabel metal4 326380 114830 331160 115196 0 FreeSans 1600 0 0 0 vddio
port 615 nsew
flabel metal4 336359 114830 341139 115196 0 FreeSans 1600 0 0 0 vddio
port 615 nsew
flabel metal4 468380 114774 473160 115224 0 FreeSans 1600 0 0 0 vssio
port 616 nsew
flabel metal4 478359 114774 483139 115224 0 FreeSans 1600 0 0 0 vssio
port 616 nsew
flabel metal5 -4 102022 316 105022 0 FreeSans 1600 90 0 0 vssd0
port 617 nsew
flabel metal5 -4 107022 316 110022 0 FreeSans 1600 90 0 0 vccd0
port 618 nsew
flabel metal5 574302 107022 574622 110022 0 FreeSans 1600 90 0 0 vccd0
port 618 nsew
flabel metal5 574302 102022 574622 105022 0 FreeSans 1600 90 0 0 vssd0
port 617 nsew
flabel metal2 561792 0 561820 300 0 FreeSans 240 90 0 0 dac_refl_to_gpio1_0[1]
port 547 nsew
flabel metal2 561904 0 561932 300 0 FreeSans 240 90 0 0 dac_refl_to_gpio1_0[0]
port 548 nsew
flabel metal2 557312 -20 557340 280 0 FreeSans 240 90 0 0 right_instramp_p_to_sio0
port 619 nsew
flabel metal2 22592 0 22620 300 0 FreeSans 240 90 0 0 adc1_comp_out
port 148 nsew
flabel metal2 22704 0 22732 300 0 FreeSans 240 90 0 0 adc1_hold
port 149 nsew
flabel metal2 22816 0 22844 300 0 FreeSans 240 90 0 0 adc1_reset
port 150 nsew
flabel metal2 22928 0 22956 300 0 FreeSans 240 90 0 0 tempsense_ena
port 151 nsew
flabel metal2 23040 0 23068 300 0 FreeSans 240 90 0 0 rdac0_ena
port 152 nsew
flabel metal2 23152 0 23180 300 0 FreeSans 240 90 0 0 rdac0_value[11]
port 153 nsew
flabel metal2 23264 0 23292 300 0 FreeSans 240 90 0 0 rdac0_value[10]
port 154 nsew
flabel metal2 23376 0 23404 300 0 FreeSans 240 90 0 0 rdac0_value[9]
port 155 nsew
flabel metal2 23488 0 23516 300 0 FreeSans 240 90 0 0 rdac0_value[8]
port 156 nsew
flabel metal2 23600 0 23628 300 0 FreeSans 240 90 0 0 rdac0_value[7]
port 157 nsew
flabel metal2 23712 0 23740 300 0 FreeSans 240 90 0 0 rdac0_value[6]
port 158 nsew
flabel metal2 23824 0 23852 300 0 FreeSans 240 90 0 0 rdac0_value[5]
port 159 nsew
flabel metal2 23936 0 23964 300 0 FreeSans 240 90 0 0 rdac0_value[4]
port 160 nsew
flabel metal2 24048 0 24076 300 0 FreeSans 240 90 0 0 rdac0_value[3]
port 161 nsew
flabel metal2 24160 0 24188 300 0 FreeSans 240 90 0 0 rdac0_value[2]
port 162 nsew
flabel metal2 24272 0 24300 300 0 FreeSans 240 90 0 0 rdac0_value[1]
port 163 nsew
flabel metal2 24384 0 24412 300 0 FreeSans 240 90 0 0 rdac0_value[0]
port 164 nsew
flabel metal2 24496 0 24524 300 0 FreeSans 240 90 0 0 rdac1_ena
port 165 nsew
flabel metal2 24608 0 24636 300 0 FreeSans 240 90 0 0 rdac1_value[11]
port 166 nsew
flabel metal2 24720 0 24748 300 0 FreeSans 240 90 0 0 rdac1_value[10]
port 167 nsew
flabel metal2 24832 0 24860 300 0 FreeSans 240 90 0 0 rdac1_value[9]
port 168 nsew
flabel metal2 24944 0 24972 300 0 FreeSans 240 90 0 0 rdac1_value[8]
port 169 nsew
flabel metal2 25056 0 25084 300 0 FreeSans 240 90 0 0 rdac1_value[7]
port 170 nsew
flabel metal2 25168 0 25196 300 0 FreeSans 240 90 0 0 rdac1_value[6]
port 171 nsew
flabel metal2 25280 0 25308 300 0 FreeSans 240 90 0 0 rdac1_value[5]
port 172 nsew
flabel metal2 25392 0 25420 300 0 FreeSans 240 90 0 0 rdac1_value[4]
port 173 nsew
flabel metal2 25504 0 25532 300 0 FreeSans 240 90 0 0 rdac1_value[3]
port 174 nsew
flabel metal2 25616 0 25644 300 0 FreeSans 240 90 0 0 rdac1_value[2]
port 175 nsew
flabel metal2 25728 0 25756 300 0 FreeSans 240 90 0 0 rdac1_value[1]
port 176 nsew
flabel metal2 25840 0 25868 300 0 FreeSans 240 90 0 0 rdac1_value[0]
port 177 nsew
flabel metal2 25952 0 25980 300 0 FreeSans 240 90 0 0 adc0_ena
port 178 nsew
flabel metal2 26064 0 26092 300 0 FreeSans 240 90 0 0 adc1_ena
port 179 nsew
flabel metal2 26176 0 26204 300 0 FreeSans 240 90 0 0 left_instramp_ena
port 180 nsew
flabel metal2 26288 0 26316 300 0 FreeSans 240 90 0 0 left_instramp_G1[4]
port 181 nsew
flabel metal2 26400 0 26428 300 0 FreeSans 240 90 0 0 left_instramp_G1[3]
port 182 nsew
flabel metal2 26512 0 26540 300 0 FreeSans 240 90 0 0 left_instramp_G1[2]
port 183 nsew
flabel metal2 26624 0 26652 300 0 FreeSans 240 90 0 0 left_instramp_G1[1]
port 184 nsew
flabel metal2 26736 0 26764 300 0 FreeSans 240 90 0 0 left_instramp_G1[0]
port 185 nsew
flabel metal2 26848 0 26876 300 0 FreeSans 240 90 0 0 left_instramp_G2[4]
port 186 nsew
flabel metal2 26960 0 26988 300 0 FreeSans 240 90 0 0 left_instramp_G2[3]
port 187 nsew
flabel metal2 27072 0 27100 300 0 FreeSans 240 90 0 0 left_instramp_G2[2]
port 188 nsew
flabel metal2 27184 0 27212 300 0 FreeSans 240 90 0 0 left_instramp_G2[1]
port 189 nsew
flabel metal2 27296 0 27324 300 0 FreeSans 240 90 0 0 left_instramp_G2[0]
port 190 nsew
flabel metal2 27408 0 27436 300 0 FreeSans 240 90 0 0 left_hgbw_opamp_ena
port 191 nsew
flabel metal2 27520 0 27548 300 0 FreeSans 240 90 0 0 left_lp_opamp_ena
port 192 nsew
flabel metal2 27632 0 27660 300 0 FreeSans 240 90 0 0 left_rheostat1_b[7]
port 193 nsew
flabel metal2 27744 0 27772 300 0 FreeSans 240 90 0 0 left_rheostat1_b[6]
port 194 nsew
flabel metal2 27856 0 27884 300 0 FreeSans 240 90 0 0 left_rheostat1_b[5]
port 195 nsew
flabel metal2 27968 0 27996 300 0 FreeSans 240 90 0 0 left_rheostat1_b[4]
port 196 nsew
flabel metal2 28080 0 28108 300 0 FreeSans 240 90 0 0 left_rheostat1_b[3]
port 197 nsew
flabel metal2 28192 0 28220 300 0 FreeSans 240 90 0 0 left_rheostat1_b[2]
port 198 nsew
flabel metal2 28304 0 28332 300 0 FreeSans 240 90 0 0 left_rheostat1_b[1]
port 199 nsew
flabel metal2 28416 0 28444 300 0 FreeSans 240 90 0 0 left_rheostat1_b[0]
port 200 nsew
flabel metal2 28528 0 28556 300 0 FreeSans 240 90 0 0 left_rheostat2_b[7]
port 201 nsew
flabel metal2 28640 0 28668 300 0 FreeSans 240 90 0 0 left_rheostat2_b[6]
port 202 nsew
flabel metal2 28752 0 28780 300 0 FreeSans 240 90 0 0 left_rheostat2_b[5]
port 203 nsew
flabel metal2 28864 0 28892 300 0 FreeSans 240 90 0 0 left_rheostat2_b[4]
port 204 nsew
flabel metal2 28976 0 29004 300 0 FreeSans 240 90 0 0 left_rheostat2_b[3]
port 205 nsew
flabel metal2 29088 0 29116 300 0 FreeSans 240 90 0 0 left_rheostat2_b[2]
port 206 nsew
flabel metal2 29200 0 29228 300 0 FreeSans 240 90 0 0 left_rheostat2_b[1]
port 207 nsew
flabel metal2 29312 0 29340 300 0 FreeSans 240 90 0 0 left_rheostat2_b[0]
port 208 nsew
flabel metal2 29424 0 29452 300 0 FreeSans 240 90 0 0 analog0_connect[1]
port 209 nsew
flabel metal2 29536 0 29564 300 0 FreeSans 240 90 0 0 analog0_connect[0]
port 210 nsew
flabel metal2 29648 0 29676 300 0 FreeSans 240 90 0 0 analog1_connect[1]
port 211 nsew
flabel metal2 29760 0 29788 276 0 FreeSans 240 90 0 0 analog1_connect[0]
port 212 nsew
flabel metal2 29872 0 29900 300 0 FreeSans 240 90 0 0 brownout_ena
port 620 nsew
flabel metal2 29984 0 30012 300 0 FreeSans 240 90 0 0 brownout_vtrip[2]
port 621 nsew
flabel metal2 30096 0 30124 300 0 FreeSans 240 90 0 0 brownout_vtrip[1]
port 622 nsew
flabel metal2 30208 0 30236 300 0 FreeSans 240 90 0 0 brownout_vtrip[0]
port 623 nsew
flabel metal2 30320 0 30348 300 0 FreeSans 240 90 0 0 brownout_otrip[2]
port 624 nsew
flabel metal2 30432 0 30460 300 0 FreeSans 240 90 0 0 brownout_otrip[1]
port 625 nsew
flabel metal2 30544 0 30572 300 0 FreeSans 240 90 0 0 brownout_otrip[0]
port 626 nsew
flabel metal2 30656 0 30684 300 0 FreeSans 240 90 0 0 brownout_isrc_sel
port 627 nsew
flabel metal2 30768 0 30796 300 0 FreeSans 240 90 0 0 brownout_oneshot
port 628 nsew
flabel metal2 30880 0 30908 300 0 FreeSans 240 90 0 0 brownout_rc_ena
port 629 nsew
flabel metal2 30992 0 31020 300 0 FreeSans 240 90 0 0 brownout_rc_dis
port 630 nsew
flabel metal2 31104 0 31132 300 0 FreeSans 240 90 0 0 brownout_vunder
port 631 nsew
flabel metal2 31216 0 31244 300 0 FreeSans 240 90 0 0 brownout_timeout
port 632 nsew
flabel metal2 31328 0 31356 300 0 FreeSans 240 90 0 0 brownout_filt
port 633 nsew
flabel metal2 31440 0 31468 300 0 FreeSans 240 90 0 0 brownout_unfilt
port 634 nsew
flabel comment s 284868 112286 284868 112286 0 FreeSans 960 90 0 0 amuxbusB_n
flabel comment s 285664 112314 285664 112314 0 FreeSans 960 90 0 0 amuxbusA_n
flabel comment s 355004 8280 355004 8280 0 FreeSans 960 90 0 0 gpio4_7_analog
flabel comment s 355526 8348 355526 8348 0 FreeSans 960 90 0 0 gpio4_6_analog
flabel comment s 356024 8368 356024 8368 0 FreeSans 960 90 0 0 gpio4_5_analog
flabel comment s 356558 8380 356558 8380 0 FreeSans 960 90 0 0 gpio4_4_analog
flabel comment s 357062 8354 357062 8354 0 FreeSans 960 90 0 0 gpio4_3_analog
flabel comment s 357592 8362 357592 8362 0 FreeSans 960 90 0 0 gpio4_2_analog
flabel comment s 358102 8374 358102 8374 0 FreeSans 960 90 0 0 gpio4_1_analog
flabel comment s 358606 8398 358606 8398 0 FreeSans 960 90 0 0 gpio4_0_analog
flabel comment s 359110 8374 359110 8374 0 FreeSans 960 90 0 0 gpio3_7_analog
flabel comment s 359632 8362 359632 8362 0 FreeSans 960 90 0 0 gpio3_6_analog
flabel comment s 360130 8398 360130 8398 0 FreeSans 960 90 0 0 gpio3_5_analog
flabel comment s 360652 8436 360652 8436 0 FreeSans 960 90 0 0 gpio3_4_analog
flabel comment s 361150 8404 361150 8404 0 FreeSans 960 90 0 0 gpio3_3_analog
flabel comment s 361684 8410 361684 8410 0 FreeSans 960 90 0 0 gpio3_2_analog
flabel comment s 362176 8424 362176 8424 0 FreeSans 960 90 0 0 gpio3_1_analog
flabel comment s 362686 8430 362686 8430 0 FreeSans 960 90 0 0 gpio3_0_analog
flabel comment s 341698 63438 341698 63438 0 FreeSans 960 0 0 0 left_vref
flabel comment s 341690 64460 341690 64460 0 FreeSans 960 0 0 0 tempsense_out
flabel comment s 341700 64976 341700 64976 0 FreeSans 960 0 0 0 dac1
flabel comment s 341688 65484 341688 65484 0 FreeSans 960 0 0 0 dac0
flabel comment s 341686 65996 341686 65996 0 FreeSans 960 0 0 0 adc1_in
flabel comment s 341676 66508 341676 66508 0 FreeSans 960 0 0 0 adc0_in
flabel comment s 341684 67020 341684 67020 0 FreeSans 960 0 0 0 comp_n
flabel comment s 341722 67532 341722 67532 0 FreeSans 960 0 0 0 comp_p
flabel comment s 341872 70092 341872 70092 0 FreeSans 960 0 0 0 left_instramp_in_n
flabel comment s 341888 70608 341888 70608 0 FreeSans 960 0 0 0 left_instramp_in_p
flabel comment s 341846 71126 341846 71126 0 FreeSans 960 0 0 0 left_lp_opamp_in_n
flabel comment s 341886 71628 341886 71628 0 FreeSans 960 0 0 0 left_lp_opamp_in_p
flabel comment s 341894 72148 341894 72148 0 FreeSans 960 0 0 0 left_hgbw_opamp_in_n
flabel comment s 341910 72654 341910 72654 0 FreeSans 960 0 0 0 left_hgbw_opamp_in_p
flabel comment s 341916 73162 341916 73162 0 FreeSans 960 0 0 0 right_hgbw_opamp_in_n
flabel comment s 341838 73680 341838 73680 0 FreeSans 960 0 0 0 right_hgbw_opamp_in_p
flabel comment s 341848 74184 341848 74184 0 FreeSans 960 0 0 0 right_lp_opamp_in_n
flabel comment s 341916 74698 341916 74698 0 FreeSans 960 0 0 0 right_lp_opamp_in_p
flabel comment s 341940 75214 341940 75214 0 FreeSans 960 0 0 0 right_instramp_in_n
flabel comment s 341522 75726 341522 75726 0 FreeSans 960 0 0 0 right_instramp_in_p
flabel comment s 571562 20800 571562 20800 0 FreeSans 960 90 0 0 vinref
flabel comment s 572196 20738 572196 20738 0 FreeSans 960 90 0 0 voutref
flabel metal3 494044 112456 494044 112456 0 FreeSans 960 0 0 0 right_instramp_out
flabel space 493978 111858 493978 111858 0 FreeSans 960 0 0 0 right_hgbw_opamp_out
flabel space 493920 111228 493920 111228 0 FreeSans 960 0 0 0 right_lp_opamp_out
flabel metal3 493910 109984 493910 109984 0 FreeSans 960 0 0 0 left_hgbw_opamp_out
flabel metal3 288992 112418 288992 112418 0 FreeSans 960 0 0 0 right_instramp_out
flabel metal3 288926 111820 288926 111820 0 FreeSans 960 0 0 0 right_hgbw_opamp_out
flabel metal3 288868 111190 288868 111190 0 FreeSans 960 0 0 0 right_lp_opamp_out
flabel metal3 288876 110568 288876 110568 0 FreeSans 960 0 0 0 left_lp_opamp_out
flabel metal3 288858 109946 288858 109946 0 FreeSans 960 0 0 0 left_hgbw_opamp_out
flabel metal3 288876 109324 288876 109324 0 FreeSans 960 0 0 0 left_instramp_out
flabel metal3 s 287234 75696 287234 75696 0 FreeSans 960 0 0 0 right_instramp_in_p
flabel metal3 s 287652 75184 287652 75184 0 FreeSans 960 0 0 0 right_instramp_in_n
flabel metal3 s 287550 73650 287550 73650 0 FreeSans 960 0 0 0 right_hgbw_opamp_in_p
flabel metal3 s 287628 73132 287628 73132 0 FreeSans 960 0 0 0 right_hgbw_opamp_in_n
flabel metal3 s 287622 72624 287622 72624 0 FreeSans 960 0 0 0 left_hgbw_opamp_in_p
flabel metal3 s 287606 72118 287606 72118 0 FreeSans 960 0 0 0 left_hgbw_opamp_in_n
flabel metal3 s 287598 71598 287598 71598 0 FreeSans 960 0 0 0 left_lp_opamp_in_p
flabel metal3 s 287558 71096 287558 71096 0 FreeSans 960 0 0 0 left_lp_opamp_in_n
flabel metal3 s 287584 70062 287584 70062 0 FreeSans 960 0 0 0 left_instramp_in_n
flabel metal3 s 287434 67502 287434 67502 0 FreeSans 960 0 0 0 comp_p
flabel metal3 s 287396 66990 287396 66990 0 FreeSans 960 0 0 0 comp_n
flabel metal3 s 287388 66478 287388 66478 0 FreeSans 960 0 0 0 adc0_in
flabel metal3 s 287398 65966 287398 65966 0 FreeSans 960 0 0 0 adc1_in
flabel metal3 s 287400 65454 287400 65454 0 FreeSans 960 0 0 0 dac0
flabel metal3 s 287412 64946 287412 64946 0 FreeSans 960 0 0 0 dac1
flabel metal3 s 287402 64430 287402 64430 0 FreeSans 960 0 0 0 tempsense_out
flabel metal3 s 287410 63408 287410 63408 0 FreeSans 960 0 0 0 left_vref
flabel metal2 5142 83610 5142 83610 0 FreeSans 960 90 0 0 adc0
flabel metal2 4542 83584 4542 83584 0 FreeSans 960 90 0 0 comp_n
flabel metal2 3942 83560 3942 83560 0 FreeSans 960 90 0 0 comp_p
flabel metal3 46514 112418 46514 112418 0 FreeSans 960 0 0 0 right_instramp_out
flabel metal3 46448 111820 46448 111820 0 FreeSans 960 0 0 0 right_hgbw_opamp_out
flabel metal3 46390 111190 46390 111190 0 FreeSans 960 0 0 0 right_lp_opamp_out
flabel metal3 46398 110568 46398 110568 0 FreeSans 960 0 0 0 left_lp_opamp_out
flabel metal3 46380 109946 46380 109946 0 FreeSans 960 0 0 0 left_hgbw_opamp_out
flabel metal3 46398 109324 46398 109324 0 FreeSans 960 0 0 0 left_instramp_out
flabel comment s 535922 75726 535922 75726 0 FreeSans 960 0 0 0 right_instramp_in_p
flabel comment s 536340 75214 536340 75214 0 FreeSans 960 0 0 0 right_instramp_in_n
flabel metal3 s 536316 74698 536316 74698 0 FreeSans 960 0 0 0 right_lp_opamp_in_p
flabel metal3 s 536248 74184 536248 74184 0 FreeSans 960 0 0 0 right_lp_opamp_in_n
flabel comment s 536238 73680 536238 73680 0 FreeSans 960 0 0 0 right_hgbw_opamp_in_p
flabel comment s 536316 73162 536316 73162 0 FreeSans 960 0 0 0 right_hgbw_opamp_in_n
flabel comment s 536310 72654 536310 72654 0 FreeSans 960 0 0 0 left_hgbw_opamp_in_p
flabel comment s 536294 72148 536294 72148 0 FreeSans 960 0 0 0 left_hgbw_opamp_in_n
flabel comment s 536286 71628 536286 71628 0 FreeSans 960 0 0 0 left_lp_opamp_in_p
flabel comment s 536246 71126 536246 71126 0 FreeSans 960 0 0 0 left_lp_opamp_in_n
flabel comment s 536288 70608 536288 70608 0 FreeSans 960 0 0 0 left_instramp_in_p
flabel comment s 536272 70092 536272 70092 0 FreeSans 960 0 0 0 left_instramp_in_n
flabel comment s 536122 67532 536122 67532 0 FreeSans 960 0 0 0 comp_p
flabel comment s 536084 67020 536084 67020 0 FreeSans 960 0 0 0 comp_n
flabel comment s 536076 66508 536076 66508 0 FreeSans 960 0 0 0 adc0_in
flabel comment s 536086 65996 536086 65996 0 FreeSans 960 0 0 0 adc1_in
flabel comment s 536106 63946 536106 63946 0 FreeSans 960 0 0 0 right_vref
flabel comment s 536098 63438 536098 63438 0 FreeSans 960 0 0 0 left_vref
flabel comment s 536102 62934 536102 62934 0 FreeSans 960 0 0 0 vinref
flabel comment s 536076 62414 536076 62414 0 FreeSans 960 0 0 0 voutref
flabel comment s 37316 74698 37316 74698 0 FreeSans 960 0 0 0 right_lp_opamp_in_p
flabel comment s 37248 74184 37248 74184 0 FreeSans 960 0 0 0 right_lp_opamp_in_n
flabel comment s 37316 73162 37316 73162 0 FreeSans 960 0 0 0 right_hgbw_opamp_in_n
flabel comment s 37310 72654 37310 72654 0 FreeSans 960 0 0 0 left_hgbw_opamp_in_p
flabel comment s 37286 71628 37286 71628 0 FreeSans 960 0 0 0 left_lp_opamp_in_p
flabel comment s 37246 71126 37246 71126 0 FreeSans 960 0 0 0 left_lp_opamp_in_n
flabel comment s 37288 70608 37288 70608 0 FreeSans 960 0 0 0 left_instramp_in_p
flabel comment s 37272 70092 37272 70092 0 FreeSans 960 0 0 0 left_instramp_in_n
flabel comment s 37122 67532 37122 67532 0 FreeSans 960 0 0 0 comp_p
flabel comment s 37084 67020 37084 67020 0 FreeSans 960 0 0 0 comp_n
flabel comment s 37076 66508 37076 66508 0 FreeSans 960 0 0 0 adc0_in
flabel comment s 37086 65996 37086 65996 0 FreeSans 960 0 0 0 adc1_in
flabel comment s 37098 63438 37098 63438 0 FreeSans 960 0 0 0 left_vref
flabel comment s 364857 18074 364857 18074 0 FreeSans 960 0 0 0 ibias50
flabel comment s 364979 16051 364979 16051 0 FreeSans 960 0 0 0 ibias100
flabel metal3 523689 9182 523689 9182 0 FreeSans 1600 0 0 0 ibias_test
flabel metal3 532128 20611 532128 20611 0 FreeSans 1600 0 0 0 vbg
flabel metal2 22256 0 22284 300 0 FreeSans 240 90 0 0 adc0_comp_out
port 144 nsew
flabel metal2 22368 0 22396 300 0 FreeSans 240 90 0 0 adc0_hold
port 145 nsew
flabel metal2 22480 0 22508 300 0 FreeSans 240 90 0 0 adc0_reset
port 146 nsew
flabel metal2 21360 0 21388 300 0 FreeSans 240 90 0 0 dac0_to_analog1
port 636 nsew
flabel metal2 21472 0 21500 300 0 FreeSans 240 90 0 0 dac1_to_analog0
port 635 nsew
flabel metal2 22144 0 22172 300 0 FreeSans 240 90 0 0 audiodac_inb
port 609 nsew
flabel metal2 22032 0 22060 300 0 FreeSans 240 90 0 0 audiodac_in
port 142 nsew
flabel metal2 21920 0 21948 300 0 FreeSans 240 90 0 0 vccd2_pwr_good
port 141 nsew
flabel metal2 21808 0 21836 300 0 FreeSans 240 90 0 0 vdda2_pwr_good
port 140 nsew
flabel metal2 21696 0 21724 300 0 FreeSans 240 90 0 0 vccd1_pwr_good
port 139 nsew
flabel metal2 21584 0 21612 300 0 FreeSans 240 90 0 0 vdda1_pwr_good
port 138 nsew
flabel metal2 21248 0 21276 300 0 FreeSans 240 90 0 0 adc1_to_analog0
port 137 nsew
flabel metal2 21136 0 21164 300 0 FreeSans 240 90 0 0 adc1_to_dac1
port 136 nsew
flabel metal2 21024 0 21052 300 0 FreeSans 240 90 0 0 adc0_to_analog1
port 135 nsew
flabel metal2 20912 0 20940 300 0 FreeSans 240 90 0 0 adc0_to_dac0
port 134 nsew
flabel metal2 20464 0 20492 300 0 FreeSans 240 90 0 0 audiodac_outb_to_analog0[1]
port 610 nsew
flabel metal2 20688 0 20716 300 0 FreeSans 240 90 0 0 audiodac_out_to_analog1[1]
port 611 nsew
flabel metal2 20576 0 20604 300 0 FreeSans 240 90 0 0 audiodac_outb_to_analog0[0]
port 667 nsew
flabel metal2 20800 0 20828 300 0 FreeSans 240 90 0 0 audiodac_out_to_analog1[0]
port 668 nsew
flabel metal2 212280 0 212308 300 0 FreeSans 240 90 0 0 adc0_dac_val[15]
port 143 nsew
flabel metal2 212168 0 212196 300 0 FreeSans 240 90 0 0 adc0_dac_val[14]
port 652 nsew
flabel metal2 212056 0 212084 300 0 FreeSans 240 90 0 0 adc0_dac_val[13]
port 653 nsew
flabel metal2 211944 0 211972 300 0 FreeSans 240 90 0 0 adc0_dac_val[12]
port 654 nsew
flabel metal2 211832 0 211860 300 0 FreeSans 240 90 0 0 adc0_dac_val[11]
port 655 nsew
flabel metal2 211720 0 211748 300 0 FreeSans 240 90 0 0 adc0_dac_val[10]
port 656 nsew
flabel metal2 211608 0 211636 300 0 FreeSans 240 90 0 0 adc0_dac_val[9]
port 657 nsew
flabel metal2 211496 0 211524 300 0 FreeSans 240 90 0 0 adc0_dac_val[8]
port 658 nsew
flabel metal2 211384 0 211412 300 0 FreeSans 240 90 0 0 adc0_dac_val[7]
port 659 nsew
flabel metal2 211272 0 211300 300 0 FreeSans 240 90 0 0 adc0_dac_val[6]
port 660 nsew
flabel metal2 211160 0 211188 300 0 FreeSans 240 90 0 0 adc0_dac_val[5]
port 661 nsew
flabel metal2 211048 0 211076 300 0 FreeSans 240 90 0 0 adc0_dac_val[4]
port 662 nsew
flabel metal2 210936 0 210964 300 0 FreeSans 240 90 0 0 adc0_dac_val[3]
port 663 nsew
flabel metal2 210824 0 210852 300 0 FreeSans 240 90 0 0 adc0_dac_val[2]
port 664 nsew
flabel metal2 210712 0 210740 300 0 FreeSans 240 90 0 0 adc0_dac_val[1]
port 665 nsew
flabel metal2 210600 0 210628 300 0 FreeSans 240 90 0 0 adc0_dac_val[0]
port 666 nsew
flabel metal2 153488 0 153516 300 0 FreeSans 240 90 0 0 adc1_dac_val[15]
port 147 nsew
flabel metal2 153376 0 153404 300 0 FreeSans 240 90 0 0 adc1_dac_val[14]
port 637 nsew
flabel metal2 153264 0 153292 300 0 FreeSans 240 90 0 0 adc1_dac_val[13]
port 638 nsew
flabel metal2 153152 0 153180 300 0 FreeSans 240 90 0 0 adc1_dac_val[12]
port 639 nsew
flabel metal2 153040 0 153068 300 0 FreeSans 240 90 0 0 adc1_dac_val[11]
port 640 nsew
flabel metal2 152928 0 152956 300 0 FreeSans 240 90 0 0 adc1_dac_val[10]
port 641 nsew
flabel metal2 152816 0 152844 300 0 FreeSans 240 90 0 0 adc1_dac_val[9]
port 642 nsew
flabel metal2 152704 0 152732 300 0 FreeSans 240 90 0 0 adc1_dac_val[8]
port 643 nsew
flabel metal2 152592 0 152620 300 0 FreeSans 240 90 0 0 adc1_dac_val[7]
port 644 nsew
flabel metal2 152480 0 152508 300 0 FreeSans 240 90 0 0 adc1_dac_val[6]
port 645 nsew
flabel metal2 152368 0 152396 300 0 FreeSans 240 90 0 0 adc1_dac_val[5]
port 646 nsew
flabel metal2 152256 0 152284 300 0 FreeSans 240 90 0 0 adc1_dac_val[4]
port 647 nsew
flabel metal2 152144 0 152172 300 0 FreeSans 240 90 0 0 adc1_dac_val[3]
port 648 nsew
flabel metal2 152032 0 152060 300 0 FreeSans 240 90 0 0 adc1_dac_val[2]
port 649 nsew
flabel metal2 151920 0 151948 300 0 FreeSans 240 90 0 0 adc1_dac_val[1]
port 650 nsew
flabel metal2 151808 0 151836 300 0 FreeSans 240 90 0 0 adc1_dac_val[0]
port 651 nsew
flabel comment s 131858 61070 131858 61070 0 FreeSans 8000 90 0 0 vccd1
flabel comment s 133148 61178 133148 61178 0 FreeSans 8000 90 0 0 vssd1
flabel comment s 131964 48228 131964 48228 0 FreeSans 8000 90 0 0 vssa1
flabel comment s 133076 48586 133076 48586 0 FreeSans 8000 90 0 0 vdda1
flabel comment s 81638 37250 81638 37250 0 FreeSans 8000 90 0 0 vssa2
flabel comment s 83108 37500 83108 37500 0 FreeSans 8000 90 0 0 vdda2
flabel metal3 528878 47843 528878 47843 0 FreeSans 1600 0 0 0 idac_snk
flabel metal3 528227 34460 528227 34460 0 FreeSans 1600 0 0 0 idac_src
flabel metal2 5726 83592 5726 83592 0 FreeSans 960 90 0 0 adc1
flabel metal2 18784 0 18812 300 0 FreeSans 240 90 0 0 left_lp_opamp_to_adc1[1]
port 119 nsew
flabel metal4 284164 102570 284164 102570 0 FreeSans 960 90 0 0 analog0_core
flabel metal4 283312 85906 283312 85906 0 FreeSans 960 90 0 0 analog1_core
flabel metal4 2928 0 3056 300 0 FreeSans 240 90 0 0 gpio6_1
port 6 nsew
flabel comment s 341786 68562 341786 68562 0 FreeSans 960 0 0 0 ulpcomp_p
flabel comment s 341758 68044 341758 68044 0 FreeSans 960 0 0 0 ulpcomp_n
flabel metal3 s 287498 68532 287498 68532 0 FreeSans 960 0 0 0 ulpcomp_p
flabel metal3 s 287470 68014 287470 68014 0 FreeSans 960 0 0 0 ulpcomp_n
flabel comment s 536186 68562 536186 68562 0 FreeSans 960 0 0 0 ulpcomp_p
flabel comment s 536158 68044 536158 68044 0 FreeSans 960 0 0 0 ulpcomp_n
flabel comment s 37158 68044 37158 68044 0 FreeSans 960 0 0 0 ulpcomp_n
flabel comment s 37186 68562 37186 68562 0 FreeSans 960 0 0 0 ulpcomp_p
flabel metal2 2766 83552 2766 83552 0 FreeSans 960 90 0 0 ulpcomp_p
flabel metal2 3358 83534 3358 83534 0 FreeSans 960 90 0 0 ulpcomp_n
flabel metal3 s 541581 5788 541581 5788 0 FreeSans 960 0 0 0 dac_vrefL
flabel metal3 s 541611 6432 541611 6432 0 FreeSans 960 0 0 0 dac_vrefH
flabel metal3 s 37268 72174 37268 72174 0 FreeSans 960 0 0 0 left_hgbw_opamp_in_n
flabel metal3 s 37212 73706 37212 73706 0 FreeSans 960 0 0 0 right_hgbw_opamp_in_p
flabel metal2 s 343106 59778 343106 59778 0 FreeSans 960 90 0 0 voutref
flabel metal2 s 343622 59762 343622 59762 0 FreeSans 960 90 0 0 vinref
flabel metal2 s 344126 59754 344126 59754 0 FreeSans 960 90 0 0 left_vref
flabel metal2 s 344632 59762 344632 59762 0 FreeSans 960 90 0 0 right_vref
flabel metal2 s 345152 59826 345152 59826 0 FreeSans 960 90 0 0 tempsense_out
flabel metal2 s 345642 59816 345642 59816 0 FreeSans 960 90 0 0 dac0
flabel metal2 s 346182 59822 346182 59822 0 FreeSans 960 90 0 0 dac1
flabel metal2 s 346696 59826 346696 59826 0 FreeSans 960 90 0 0 vbgtc
flabel metal2 s 347202 59832 347202 59832 0 FreeSans 960 90 0 0 vbgsc
flabel metal2 s 348734 59836 348734 59836 0 FreeSans 960 90 0 0 adc0_in
flabel metal2 s 349246 59848 349246 59848 0 FreeSans 960 90 0 0 adc1_in
flabel metal2 s 349766 59866 349766 59866 0 FreeSans 960 90 0 0 comp_n
flabel metal2 s 350298 59890 350298 59890 0 FreeSans 960 90 0 0 comp_p
flabel metal2 s 351282 59910 351282 59910 0 FreeSans 960 90 0 0 ulpcomp_p
flabel metal2 s 350790 59900 350790 59900 0 FreeSans 960 90 0 0 ulpcomp_n
flabel metal3 274234 19474 274234 19474 0 FreeSans 960 0 0 0 audiodac_out
flabel metal3 274220 32536 274220 32536 0 FreeSans 960 0 0 0 audiodac_outb
flabel metal3 413828 61854 413828 61854 0 FreeSans 960 0 0 0 vcmosref
flabel metal3 423992 18588 423992 18588 0 FreeSans 960 0 0 0 brownout_ibias
flabel metal3 332424 60272 332424 60272 0 FreeSans 960 0 0 0 ibias_comp
flabel metal3 456254 21226 456254 21226 0 FreeSans 960 0 0 0 left_lp_opamp_ibias
flabel metal3 456020 20796 456020 20796 0 FreeSans 960 0 0 0 right_lp_opamp_ibias
flabel metal4 388462 24166 388462 24166 0 FreeSans 960 90 0 0 left_hgbw_opamp_ibias
flabel metal4 435530 24310 435530 24310 0 FreeSans 960 90 0 0 ibias_ov
flabel space 437094 18660 437094 18660 0 FreeSans 960 0 0 0 user_ibias50
flabel metal4 434782 16216 434782 16216 0 FreeSans 960 0 0 0 user_ibias100
flabel metal3 454150 18408 454150 18408 0 FreeSans 960 90 0 0 ibias_instr1
flabel metal3 452570 18402 452570 18402 0 FreeSans 960 90 0 0 ibias_instr2
flabel metal3 417878 18262 417878 18262 0 FreeSans 960 90 0 0 ibias_idac
flabel metal4 477444 16626 477444 16626 0 FreeSans 960 0 0 0 ibias_test
flabel metal3 550596 61824 550596 61824 0 FreeSans 1280 0 0 0 sio0_core
flabel metal3 550544 61390 550544 61390 0 FreeSans 1280 0 0 0 sio1_core
flabel metal4 388888 24234 388888 24234 0 FreeSans 960 90 0 0 right_hgbw_opamp_ibias
flabel metal2 540268 0 540338 300 0 FreeSans 240 90 0 0 porb_h[1]
port 355 nsew
flabel metal2 31561 0 31631 300 0 FreeSans 240 90 0 0 porb_h[0]
port 669 nsew
flabel metal2 387420 39346 387420 39346 0 FreeSans 1600 0 0 0 vbgpwr
flabel metal4 572144 0 572272 300 0 FreeSans 240 90 0 0 gpio2_3
port 556 nsew
flabel metal4 571632 0 571760 300 0 FreeSans 240 90 0 0 gpio2_2
port 557 nsew
flabel metal4 571120 0 571248 300 0 FreeSans 240 90 0 0 gpio2_1
port 558 nsew
flabel metal4 570608 0 570736 300 0 FreeSans 240 90 0 0 gpio2_0
port 559 nsew
flabel metal4 570096 0 570224 300 0 FreeSans 240 90 0 0 gpio1_7
port 560 nsew
flabel metal4 569584 0 569712 300 0 FreeSans 240 90 0 0 gpio1_6
port 561 nsew
flabel metal4 569072 0 569200 300 0 FreeSans 240 90 0 0 gpio1_5
port 562 nsew
flabel metal4 568560 0 568688 300 0 FreeSans 240 90 0 0 gpio1_4
port 563 nsew
flabel metal4 568048 0 568176 300 0 FreeSans 240 90 0 0 right_vref
port 564 nsew
flabel metal4 567536 0 567664 300 0 FreeSans 240 90 0 0 gpio1_3
port 565 nsew
flabel metal4 567024 0 567152 300 0 FreeSans 240 90 0 0 gpio1_2
port 566 nsew
flabel metal4 566512 0 566640 300 0 FreeSans 240 90 0 0 gpio1_1
port 567 nsew
flabel metal4 566000 0 566128 300 0 FreeSans 240 90 0 0 gpio1_0
port 568 nsew
flabel comment s 570298 46786 570298 46786 0 FreeSans 960 90 0 0 right_vref
flabel metal4 80812 114900 81012 115200 0 FreeSans 480 90 0 0 gpio4_4
port 576 nsew
flabel comment s 100214 52344 100214 52344 0 FreeSans 8000 90 0 0 vccd2
flabel comment s 94180 52621 94180 52621 0 FreeSans 8000 90 0 0 vssd2
flabel metal4 503812 114900 504012 115200 0 FreeSans 480 90 0 0 gpio3_3
port 589 nsew
flabel metal3 s 287600 70578 287600 70578 0 FreeSans 960 0 0 0 left_instramp_in_p
flabel metal3 s 17309 7010 17309 7010 0 FreeSans 960 0 0 0 adc_vrefL
flabel metal3 s 17280 7638 17280 7638 0 FreeSans 960 0 0 0 adc_vrefH
flabel comment s 341713 63967 341713 63967 0 FreeSans 960 0 0 0 right_vref
flabel metal2 19792 0 19820 300 0 FreeSans 240 90 0 0 right_instramp_p_to_left_rheostat2_out
port 128 nsew
flabel metal2 552496 0 552524 300 0 FreeSans 240 90 0 0 right_instramp_p_to_right_rheostat1_out
port 464 nsew
flabel metal2 553280 0 553308 300 0 FreeSans 240 90 0 0 right_instramp_n_to_right_rheostat1_out
port 471 nsew
flabel metal2 17664 0 17692 300 0 FreeSans 240 90 0 0 left_instramp_p_to_left_rheostat1_out
port 109 nsew
flabel metal2 18112 0 18140 300 0 FreeSans 240 90 0 0 left_instramp_n_to_left_rheostat1_out
port 113 nsew
flabel metal2 20240 0 20268 300 0 FreeSans 240 90 0 0 right_instramp_n_to_left_rheostat2_out
port 132 nsew
flabel metal2 551040 0 551068 300 0 FreeSans 240 90 0 0 left_instramp_n_to_right_rheostat2_out
port 451 nsew
flabel metal2 550144 0 550172 300 0 FreeSans 240 90 0 0 left_instramp_p_to_right_rheostat2_out
port 443 nsew
<< properties >>
string FIXED_BBOX 0 0 574978 115318
<< end >>
