** sch_path: /home/tim/gits/frigate_analog/xschem/frigate_analog.sch
.subckt frigate_analog left_hgbw_opamp_p_to_gpio5_2[1] left_hgbw_opamp_p_to_gpio5_2[0] ibias_test_to_gpio1_2[1]
+ ibias_test_to_gpio1_2[0] right_lp_opamp_p_to_dac0 overvoltage_ena left_instramp_to_ulpcomp_p[1] left_instramp_to_ulpcomp_p[0] vdda0
+ right_lp_opamp_p_to_analog0 vssa0 left_hgbw_opamp_p_to_dac0 left_instramp_to_comp_p[1] left_instramp_to_comp_p[0] overvoltage_trim[3] overvoltage_trim[2]
+ overvoltage_trim[1] overvoltage_trim[0] vbg_test_to_gpio1_1[1] vbg_test_to_gpio1_1[0] vdda1 overvoltage_out left_instramp_to_adc0[1]
+ left_instramp_to_adc0[0] right_lp_opamp_p_to_amuxbusA left_hgbw_opamp_p_to_analog0 idac_to_gpio1_3[1] idac_to_gpio1_3[0]
+ left_instramp_p_to_left_rheostat1_out left_hgbw_opamp_p_to_amuxbusA vssa1 tempsense_ena left_instramp_to_gpio4_4[1] left_instramp_to_gpio4_4[0] idac_to_gpio1_2[1]
+ idac_to_gpio1_2[0] vdda2 left_instramp_to_analog1[1] left_instramp_to_analog1[0] left_instramp_p_to_right_rheostat2_out right_lp_opamp_p_to_sio0
+ adc_refh_to_gpio6_6[1] adc_refh_to_gpio6_6[0] vdda1_pwr_good left_hgbw_opamp_p_to_sio0 left_instramp_to_amuxbusB[1] left_instramp_to_amuxbusB[0]
+ right_lp_opamp_p_to_tempsense vssa2 dac_refh_to_gpio1_1[1] dac_refh_to_gpio1_1[0] vccd1_pwr_good right_instramp_to_ulpcomp_n[1] right_instramp_to_ulpcomp_n[0]
+ left_hgbw_opamp_p_to_left_vref vccd1 right_lp_opamp_p_to_left_vref adc_refl_to_gpio6_7[1] adc_refl_to_gpio6_7[0] vdda2_pwr_good right_lp_opamp_p_to_voutref
+ vssd1 left_hgbw_opamp_p_to_voutref right_instramp_to_comp_n[1] right_instramp_to_comp_n[0] dac_refl_to_gpio1_0[1]
+ dac_refl_to_gpio1_0[0] vccd2_pwr_good right_lp_opamp_p_to_gpio2_5[1] right_lp_opamp_p_to_gpio2_5[0] right_instramp_to_adc1[1] right_instramp_to_adc1[0]
+ left_hgbw_opamp_p_to_gpio2_1[1] left_hgbw_opamp_p_to_gpio2_1[0] vccd2 right_lp_opamp_to_ulpcomp_p[1] right_lp_opamp_to_ulpcomp_p[0] right_lp_opamp_n_to_dac1
+ right_instramp_to_analog0[1] right_instramp_to_analog0[0] vssd2 left_hgbw_opamp_n_to_gpio5_3[1] left_hgbw_opamp_n_to_gpio5_3[0] right_lp_opamp_to_comp_p[1]
+ right_lp_opamp_to_comp_p[0] right_instramp_to_amuxbusA[1] right_instramp_to_amuxbusA[0] right_lp_opamp_n_to_analog1 left_hgbw_opamp_n_to_dac1
+ right_lp_opamp_to_adc0[1] right_lp_opamp_to_adc0[0] right_lp_opamp_n_to_amuxbusB left_hgbw_opamp_n_to_analog1 right_instramp_to_gpio3_0[1]
+ right_instramp_to_gpio3_0[0] right_lp_opamp_to_gpio4_7[1] right_lp_opamp_to_gpio4_7[0] left_instramp_n_to_gpio5_7[1] left_instramp_n_to_gpio5_7[0]
+ right_instramp_n_to_left_rheostat2_out left_hgbw_opamp_n_to_amuxbusB idac_value[11] idac_value[10] idac_value[9] idac_value[8] idac_value[7] idac_value[6] idac_value[5]
+ idac_value[4] idac_value[3] idac_value[2] idac_value[1] idac_value[0] right_lp_opamp_to_gpio4_3[1] right_lp_opamp_to_gpio4_3[0]
+ left_instramp_ena right_lp_opamp_n_to_rheostat_tap left_instramp_n_to_analog1 left_instramp_n_to_right_rheostat2_out right_lp_opamp_to_analog1[1]
+ right_lp_opamp_to_analog1[0] idac_ena left_instramp_G1[4] left_instramp_G1[3] left_instramp_G1[2] left_instramp_G1[1] left_instramp_G1[0]
+ left_hgbw_opamp_n_to_rheostat_tap right_lp_opamp_n_to_sio1 left_instramp_n_to_amuxbusB right_lp_opamp_to_amuxbusB[1] right_lp_opamp_to_amuxbusB[0] audiodac_in
+ left_instramp_G2[4] left_instramp_G2[3] left_instramp_G2[2] left_instramp_G2[1] left_instramp_G2[0] right_lp_opamp_n_to_vbgtc left_instramp_n_to_sio1
+ left_hgbw_opamp_n_to_sio1 right_lp_opamp_to_gpio3_7[1] right_lp_opamp_to_gpio3_7[0] rdac0_ena left_hgbw_opamp_ena left_hgbw_opamp_n_to_vbgtc
+ left_instramp_n_to_right_vref right_lp_opamp_n_to_right_vref right_lp_opamp_to_gpio3_3[1] right_lp_opamp_to_gpio3_3[0] rdac0_value[11] rdac0_value[10]
+ rdac0_value[9] rdac0_value[8] rdac0_value[7] rdac0_value[6] rdac0_value[5] rdac0_value[4] rdac0_value[3] rdac0_value[2] rdac0_value[1]
+ rdac0_value[0] left_lp_opamp_ena left_hgbw_opamp_n_to_right_vref left_instramp_n_to_vinref right_lp_opamp_n_to_vinref
+ right_hgbw_opamp_to_ulpcomp_n[1] right_hgbw_opamp_to_ulpcomp_n[0] rdac1_ena left_rheostat1_b[7] left_rheostat1_b[6] left_rheostat1_b[5] left_rheostat1_b[4]
+ left_rheostat1_b[3] left_rheostat1_b[2] left_rheostat1_b[1] left_rheostat1_b[0] right_lp_opamp_n_to_gpio2_4[1] right_lp_opamp_n_to_gpio2_4[0]
+ left_hgbw_opamp_n_to_vinref rdac1_value[11] rdac1_value[10] rdac1_value[9] rdac1_value[8] rdac1_value[7] rdac1_value[6] rdac1_value[5] rdac1_value[4]
+ rdac1_value[3] rdac1_value[2] rdac1_value[1] rdac1_value[0] right_hgbw_opamp_to_comp_n[1] right_hgbw_opamp_to_comp_n[0] left_rheostat2_b[7]
+ left_rheostat2_b[6] left_rheostat2_b[5] left_rheostat2_b[4] left_rheostat2_b[3] left_rheostat2_b[2] left_rheostat2_b[1] left_rheostat2_b[0]
+ left_instramp_p_to_gpio5_6[1] left_instramp_p_to_gpio5_6[0] left_hgbw_opamp_n_to_gpio2_0[1] left_hgbw_opamp_n_to_gpio2_0[0] right_hgbw_opamp_p_to_gpio5_0[1]
+ right_hgbw_opamp_p_to_gpio5_0[0] right_hgbw_opamp_to_adc1[1] right_hgbw_opamp_to_adc1[0] adc0_ena left_lp_opamp_p_to_dac0 left_instramp_p_to_analog0
+ right_instramp_ena right_hgbw_opamp_p_to_dac0 right_hgbw_opamp_to_gpio4_6[1] right_hgbw_opamp_to_gpio4_6[0] adc0_reset left_instramp_p_to_amuxbusA
+ left_lp_opamp_p_to_analog0 right_instramp_G1[4] right_instramp_G1[3] right_instramp_G1[2] right_instramp_G1[1] right_instramp_G1[0]
+ right_hgbw_opamp_p_to_analog0 right_hgbw_opamp_to_gpio4_2[1] right_hgbw_opamp_to_gpio4_2[0] adc0_hold right_hgbw_opamp_p_to_amuxbusA left_instramp_p_to_sio0
+ right_instramp_G2[4] right_instramp_G2[3] right_instramp_G2[2] right_instramp_G2[1] right_instramp_G2[0] left_lp_opamp_p_to_amuxbusA
+ right_hgbw_opamp_to_analog0[1] right_hgbw_opamp_to_analog0[0] adc0_dac_val[15] adc0_dac_val[14] adc0_dac_val[13] adc0_dac_val[12] adc0_dac_val[11]
+ adc0_dac_val[10] adc0_dac_val[9] adc0_dac_val[8] adc0_dac_val[7] adc0_dac_val[6] adc0_dac_val[5] adc0_dac_val[4] adc0_dac_val[3] adc0_dac_val[2]
+ adc0_dac_val[1] adc0_dac_val[0] left_instramp_p_to_tempsense right_instramp_p_to_left_rheostat2_out right_hgbw_opamp_ena
+ right_instramp_p_to_right_rheostat1_out right_hgbw_opamp_to_amuxbusA[1] right_hgbw_opamp_to_amuxbusA[0] adc0_comp_out left_instramp_p_to_left_vref right_lp_opamp_ena
+ left_lp_opamp_p_to_sio0 right_hgbw_opamp_p_to_sio0 right_hgbw_opamp_to_gpio3_6[1] right_hgbw_opamp_to_gpio3_6[0] adc1_ena left_hgbw_opamp_p_to_tempsense
+ right_rheostat1_b[7] right_rheostat1_b[6] right_rheostat1_b[5] right_rheostat1_b[4] right_rheostat1_b[3] right_rheostat1_b[2] right_rheostat1_b[1]
+ right_rheostat1_b[0] left_instramp_p_to_voutref right_hgbw_opamp_p_to_left_vref right_hgbw_opamp_to_gpio3_2[1] right_hgbw_opamp_to_gpio3_2[0]
+ adc1_reset right_instramp_n_to_analog1 right_rheostat2_b[7] right_rheostat2_b[6] right_rheostat2_b[5] right_rheostat2_b[4]
+ right_rheostat2_b[3] right_rheostat2_b[2] right_rheostat2_b[1] right_rheostat2_b[0] left_lp_opamp_p_to_left_vref right_hgbw_opamp_p_to_voutref
+ left_hgbw_opamp_to_ulpcomp_p[1] left_hgbw_opamp_to_ulpcomp_p[0] right_instramp_n_to_amuxbusB left_lp_opamp_p_to_voutref right_hgbw_opamp_p_to_gpio2_3[1]
+ right_hgbw_opamp_p_to_gpio2_3[0] adc1_hold left_hgbw_opamp_to_comp_p[1] left_hgbw_opamp_to_comp_p[0] left_lp_opamp_n_to_gpio5_5[1] left_lp_opamp_n_to_gpio5_5[0]
+ right_instramp_n_to_sio1 right_hgbw_opamp_n_to_gpio5_1[1] right_hgbw_opamp_n_to_gpio5_1[0] adc1_dac_val[15] adc1_dac_val[14] adc1_dac_val[13]
+ adc1_dac_val[12] adc1_dac_val[11] adc1_dac_val[10] adc1_dac_val[9] adc1_dac_val[8] adc1_dac_val[7] adc1_dac_val[6] adc1_dac_val[5] adc1_dac_val[4]
+ adc1_dac_val[3] adc1_dac_val[2] adc1_dac_val[1] adc1_dac_val[0] left_hgbw_opamp_to_adc0[1] left_hgbw_opamp_to_adc0[0]
+ right_instramp_n_to_right_vref comp_ena left_lp_opamp_n_to_dac1 adc1_comp_out right_hgbw_opamp_n_to_dac1 left_hgbw_opamp_to_gpio4_5[1]
+ left_hgbw_opamp_to_gpio4_5[0] comp_trim[5] comp_trim[4] comp_trim[3] comp_trim[2] comp_trim[1] comp_trim[0] right_instramp_n_to_vinref
+ left_lp_opamp_n_to_analog1 right_hgbw_opamp_n_to_analog1 left_hgbw_opamp_to_gpio4_1[1] left_hgbw_opamp_to_gpio4_1[0] left_lp_opamp_n_to_amuxbusB
+ comp_hyst[1] comp_hyst[0] right_instramp_n_to_gpio2_6[1] right_instramp_n_to_gpio2_6[0] right_hgbw_opamp_n_to_amuxbusB
+ left_hgbw_opamp_to_analog1[1] left_hgbw_opamp_to_analog1[0] comp_out right_instramp_p_to_analog0 left_instramp_n_to_left_rheostat1_out
+ right_instramp_n_to_right_rheostat1_out left_hgbw_opamp_to_amuxbusB[1] left_hgbw_opamp_to_amuxbusB[0] ulpcomp_ena right_instramp_p_to_amuxbusA
+ right_hgbw_opamp_n_to_rheostat_tap left_lp_opamp_n_to_rheostat_tap left_hgbw_opamp_to_gpio3_5[1] left_hgbw_opamp_to_gpio3_5[0] right_instramp_p_to_tempsense
+ ulpcomp_clk left_lp_opamp_n_to_sio1 right_hgbw_opamp_n_to_sio1 left_hgbw_opamp_to_gpio3_1[1] left_hgbw_opamp_to_gpio3_1[0]
+ right_instramp_p_to_left_vref left_lp_opamp_n_to_vbgsc right_hgbw_opamp_n_to_vbgsc ulpcomp_out left_lp_opamp_to_ulpcomp_n[1] left_lp_opamp_to_ulpcomp_n[0]
+ right_instramp_p_to_voutref left_lp_opamp_n_to_right_vref right_hgbw_opamp_n_to_right_vref left_lp_opamp_to_comp_n[1] left_lp_opamp_to_comp_n[0]
+ right_instramp_p_to_gpio2_7[1] right_instramp_p_to_gpio2_7[0] left_lp_opamp_n_to_vinref right_hgbw_opamp_n_to_vinref left_lp_opamp_to_adc1[1]
+ left_lp_opamp_to_adc1[0] left_lp_opamp_p_to_gpio5_4[1] left_lp_opamp_p_to_gpio5_4[0] right_hgbw_opamp_n_to_gpio2_2[1] right_hgbw_opamp_n_to_gpio2_2[0]
+ bandgap_ena bandgap_trim[15] bandgap_trim[14] bandgap_trim[13] bandgap_trim[12] bandgap_trim[11] bandgap_trim[10] bandgap_trim[9]
+ bandgap_trim[8] bandgap_trim[7] bandgap_trim[6] bandgap_trim[5] bandgap_trim[4] bandgap_trim[3] bandgap_trim[2] bandgap_trim[1] bandgap_trim[0]
+ left_lp_opamp_to_gpio4_0[1] left_lp_opamp_to_gpio4_0[0] ldo_ena left_lp_opamp_to_analog0[1] left_lp_opamp_to_analog0[0] ibias_ena
+ left_lp_opamp_to_amuxbusA[1] left_lp_opamp_to_amuxbusA[0] ibias_src_ena[23] ibias_src_ena[22] ibias_src_ena[21] ibias_src_ena[20] ibias_src_ena[19]
+ ibias_src_ena[18] ibias_src_ena[17] ibias_src_ena[16] ibias_src_ena[15] ibias_src_ena[14] ibias_src_ena[13] ibias_src_ena[12] ibias_src_ena[11]
+ ibias_src_ena[10] ibias_src_ena[9] ibias_src_ena[8] ibias_src_ena[7] ibias_src_ena[6] ibias_src_ena[5] ibias_src_ena[4] ibias_src_ena[3]
+ ibias_src_ena[2] ibias_src_ena[1] ibias_src_ena[0] left_lp_opamp_to_gpio3_4[1] left_lp_opamp_to_gpio3_4[0] ibias_snk_ena[3] ibias_snk_ena[2]
+ ibias_snk_ena[1] ibias_snk_ena[0] ibias_ref_select por porb porb_h[1] porb_h[0] gpio1_0 user_voutref gpio4_0 ulpcomp_p_to_dac0 adc0_to_dac0
+ gpio4_1 gpio1_1 user_vinref ulpcomp_p_to_analog1 adc0_to_analog1 gpio4_2 user_left_vref gpio1_2 ulpcomp_p_to_sio0 adc0_to_vbgtc gpio4_3
+ gpio1_3 user_right_vref ulpcomp_p_to_vbgtc adc0_to_tempsense gpio1_4 gpio4_4 user_tempsense ulpcomp_p_to_tempsense adc0_to_left_vref
+ gpio4_5 gpio1_5 user_dac0 ulpcomp_p_to_left_vref adc0_to_voutref gpio4_6 gpio1_6 user_dac1 ulpcomp_p_to_voutref adc0_to_gpio6_4[1]
+ adc0_to_gpio6_4[0] gpio4_7 gpio1_7 user_vbgtc ulpcomp_p_to_gpio6_0[1] ulpcomp_p_to_gpio6_0[0] adc0_to_gpio1_3[1] adc0_to_gpio1_3[0] gpio5_0 gpio2_0
+ user_vbgsc ulpcomp_p_to_gpio1_7[1] ulpcomp_p_to_gpio1_7[0] adc1_to_dac1 user_ibias50 gpio5_1 gpio2_1 ulpcomp_n_to_dac1 adc1_to_analog0
+ user_ibias100 gpio5_2 gpio2_2 ulpcomp_n_to_analog0 adc1_to_vbgsc gpio5_3 gpio2_3 user_adc0 ulpcomp_n_to_sio1 adc1_to_right_vref gpio2_4 gpio5_4
+ user_adc1 ulpcomp_n_to_vbgsc adc1_to_vinref gpio5_5 gpio2_5 user_comp_n ulpcomp_n_to_right_vref adc1_to_gpio6_5[1] adc1_to_gpio6_5[0]
+ gpio5_6 gpio2_6 user_comp_p ulpcomp_n_to_vinref adc1_to_gpio1_2[1] adc1_to_gpio1_2[0] gpio5_7 gpio2_7 user_ulpcomp_n
+ ulpcomp_n_to_gpio6_1[1] ulpcomp_n_to_gpio6_1[0] sio0_connect[1] sio0_connect[0] gpio6_0 gpio3_0 user_ulpcomp_p ulpcomp_n_to_gpio1_6[1]
+ ulpcomp_n_to_gpio1_6[0] sio1_connect[1] sio1_connect[0] gpio6_1 gpio3_1 comp_p_to_dac0 user_gpio3_0_analog analog0_connect[1] analog0_connect[0] gpio6_2
+ gpio3_2 comp_p_to_analog1 user_gpio3_1_analog analog1_connect[1] analog1_connect[0] gpio6_3 gpio3_3 comp_p_to_sio0 user_gpio3_2_analog
+ vbgtc_to_user gpio3_4 gpio6_4 comp_p_to_vbgtc user_gpio3_3_analog vbgsc_to_user gpio6_5 gpio3_5 comp_p_to_tempsense user_gpio3_4_analog
+ user_to_comp_n[1] user_to_comp_n[0] gpio6_6 gpio3_6 comp_p_to_left_vref user_gpio3_5_analog user_to_comp_p[1] user_to_comp_p[0] gpio6_7 gpio3_7
+ comp_p_to_voutref user_gpio3_6_analog user_to_ulpcomp_n[1] user_to_ulpcomp_n[0] analog0 sio0 comp_p_to_gpio6_2[1] comp_p_to_gpio6_2[0]
+ user_gpio3_7_analog user_to_ulpcomp_p[1] user_to_ulpcomp_p[0] analog1 sio1 comp_p_to_gpio1_5[1] comp_p_to_gpio1_5[0] user_gpio4_0_analog
+ user_to_adc0[1] user_to_adc0[0] comp_n_to_dac1 user_gpio4_1_analog user_to_adc1[1] user_to_adc1[0] comp_n_to_analog0 user_gpio4_2_analog
+ dac0_to_user voutref user_gpio4_3_analog dac1_to_user vbg comp_n_to_sio1 ibias_lsxo vinref user_gpio4_4_analog tempsense_to_user
+ comp_n_to_vbgsc ibias_hsxo right_vref user_gpio4_5_analog right_vref_to_user comp_n_to_right_vref left_vref user_gpio4_6_analog left_vref_to_user
+ comp_n_to_vinref user_gpio4_7_analog vinref_to_user comp_n_to_gpio6_3[1] comp_n_to_gpio6_3[0] voutref_to_user comp_n_to_gpio1_4[1]
+ comp_n_to_gpio1_4[0] right_instramp_p_to_sio0 dac0_to_analog1 dac1_to_analog0 audiodac_out_to_analog1[1] audiodac_out_to_analog1[0]
+ audiodac_outb_to_analog0[1] audiodac_outb_to_analog0[0] audiodac_inb vddio vssio tempsense_sel ldo_ref_sel bandgap_sel brownout_vunder brownout_timeout
+ brownout_filt brownout_unfilt brownout_ena brownout_vtrip[2] brownout_vtrip[1] brownout_vtrip[0] brownout_otrip[2] brownout_otrip[1]
+ brownout_otrip[0] brownout_isrc_sel brownout_oneshot brownout_rc_ena brownout_rc_dis amuxbus_a_n amuxbus_b_n vccd0 vssd0
*.PININFO vdda0:B left_instramp_ena:I vssa0:B vdda1:B vssa1:B vdda2:B vssa2:B vccd1:B vssd1:B vccd2:B vssd2:B
*+ left_instramp_G1[4:0]:I left_instramp_G2[4:0]:I left_hgbw_opamp_ena:I left_lp_opamp_ena:I left_rheostat1_b[7:0]:I left_rheostat2_b[7:0]:I
*+ right_instramp_ena:I right_instramp_G1[4:0]:I right_instramp_G2[4:0]:I right_hgbw_opamp_ena:I right_lp_opamp_ena:I right_rheostat1_b[7:0]:I
*+ right_rheostat2_b[7:0]:I comp_ena:I comp_trim[5:0]:I comp_hyst[1:0]:I comp_out:O ulpcomp_ena:I ulpcomp_out:O ulpcomp_clk:I bandgap_ena:I
*+ bandgap_trim[15:0]:I ldo_ena:I ibias_ena:I ibias_src_ena[23:0]:I ibias_snk_ena[3:0]:I ibias_ref_select:I por:O porb:O porb_h[1:0]:O overvoltage_ena:I
*+ overvoltage_trim[3:0]:I overvoltage_out:O tempsense_ena:I vdda1_pwr_good:O vccd1_pwr_good:O vdda2_pwr_good:O vccd2_pwr_good:O idac_value[11:0]:I
*+ idac_ena:I audiodac_in:I rdac0_ena:I rdac0_value[11:0]:I rdac1_ena:I rdac1_value[11:0]:I adc0_ena:I adc0_reset:I adc0_hold:I
*+ adc0_dac_val[15:0]:I adc0_comp_out:O adc1_ena:I adc1_reset:I adc1_hold:I adc1_dac_val[15:0]:I adc1_comp_out:O ibias_test_to_gpio1_2[1:0]:I
*+ vbg_test_to_gpio1_1[1:0]:I idac_to_gpio1_3[1:0]:I idac_to_gpio1_2[1:0]:I adc_refh_to_gpio6_6[1:0]:I dac_refh_to_gpio1_1[1:0]:I adc_refl_to_gpio6_7[1:0]:I
*+ dac_refl_to_gpio1_0[1:0]:I right_lp_opamp_to_ulpcomp_p[1:0]:I right_lp_opamp_to_comp_p[1:0]:I right_lp_opamp_to_adc0[1:0]:I right_lp_opamp_to_gpio4_7[1:0]:I
*+ right_lp_opamp_to_analog1[1:0]:I right_lp_opamp_to_amuxbusB[1:0]:I right_lp_opamp_to_gpio3_7[1:0]:I right_lp_opamp_to_gpio3_3[1:0]:I
*+ right_lp_opamp_to_gpio4_3[1:0]:I right_hgbw_opamp_to_ulpcomp_n[1:0]:I right_hgbw_opamp_to_comp_n[1:0]:I right_hgbw_opamp_to_adc1[1:0]:I
*+ right_hgbw_opamp_to_gpio4_6[1:0]:I right_hgbw_opamp_to_analog0[1:0]:I right_hgbw_opamp_to_amuxbusA[1:0]:I right_hgbw_opamp_to_gpio3_6[1:0]:I
*+ right_hgbw_opamp_to_gpio3_2[1:0]:I right_hgbw_opamp_to_gpio4_2[1:0]:I left_hgbw_opamp_to_ulpcomp_p[1:0]:I left_hgbw_opamp_to_comp_p[1:0]:I
*+ left_hgbw_opamp_to_adc0[1:0]:I left_hgbw_opamp_to_gpio4_5[1:0]:I left_hgbw_opamp_to_analog1[1:0]:I left_hgbw_opamp_to_amuxbusB[1:0]:I
*+ left_hgbw_opamp_to_gpio3_5[1:0]:I left_hgbw_opamp_to_gpio3_1[1:0]:I left_hgbw_opamp_to_gpio4_1[1:0]:I left_lp_opamp_to_ulpcomp_n[1:0]:I
*+ left_lp_opamp_to_comp_n[1:0]:I left_lp_opamp_to_adc1[1:0]:I left_lp_opamp_to_analog0[1:0]:I left_lp_opamp_to_amuxbusA[1:0]:I left_lp_opamp_to_gpio3_4[1:0]:I
*+ left_lp_opamp_to_gpio4_0[1:0]:I right_lp_opamp_p_to_dac0:I right_lp_opamp_p_to_analog0:I right_lp_opamp_p_to_amuxbusA:I left_instramp_p_to_left_rheostat1_out:I
*+ right_lp_opamp_p_to_tempsense:I right_lp_opamp_p_to_left_vref:I right_lp_opamp_p_to_voutref:I right_lp_opamp_p_to_gpio2_5[1:0]:I right_lp_opamp_p_to_sio0:I
*+ right_lp_opamp_n_to_dac1:I right_lp_opamp_n_to_analog1:I right_lp_opamp_n_to_amuxbusB:I right_instramp_n_to_left_rheostat2_out:I right_lp_opamp_n_to_vbgtc:I
*+ right_lp_opamp_n_to_right_vref:I right_lp_opamp_n_to_vinref:I right_lp_opamp_n_to_gpio2_4[1:0]:I right_lp_opamp_n_to_sio1:I right_hgbw_opamp_p_to_dac0:I
*+ right_hgbw_opamp_p_to_analog0:I right_hgbw_opamp_p_to_amuxbusA:I right_instramp_p_to_right_rheostat1_out:I right_hgbw_opamp_p_to_left_vref:I
*+ right_hgbw_opamp_p_to_voutref:I right_hgbw_opamp_p_to_gpio2_3[1:0]:I right_hgbw_opamp_p_to_sio0:I right_lp_opamp_n_to_rheostat_tap:I
*+ right_hgbw_opamp_p_to_gpio5_0[1:0]:I right_hgbw_opamp_n_to_dac1:I right_hgbw_opamp_n_to_analog1:I right_hgbw_opamp_n_to_amuxbusB:I
*+ right_instramp_n_to_right_rheostat1_out:I right_hgbw_opamp_n_to_vbgsc:I right_hgbw_opamp_n_to_right_vref:I right_hgbw_opamp_n_to_vinref:I
*+ right_hgbw_opamp_n_to_gpio2_2[1:0]:I right_hgbw_opamp_n_to_sio1:I right_hgbw_opamp_n_to_rheostat_tap:I right_hgbw_opamp_n_to_gpio5_1[1:0]:I
*+ left_hgbw_opamp_p_to_gpio5_2[1:0]:I left_hgbw_opamp_p_to_dac0:I left_hgbw_opamp_p_to_analog0:I left_hgbw_opamp_p_to_amuxbusA:I
*+ left_instramp_p_to_right_rheostat2_out:I left_hgbw_opamp_p_to_sio0:I left_hgbw_opamp_p_to_tempsense:I left_hgbw_opamp_p_to_left_vref:I left_hgbw_opamp_p_to_voutref:I
*+ left_hgbw_opamp_p_to_gpio2_1[1:0]:I left_hgbw_opamp_n_to_gpio5_3[1:0]:I left_hgbw_opamp_n_to_dac1:I left_hgbw_opamp_n_to_analog1:I left_hgbw_opamp_n_to_amuxbusB:I
*+ left_instramp_n_to_right_rheostat2_out:I left_hgbw_opamp_n_to_rheostat_tap:I left_hgbw_opamp_n_to_sio1:I left_hgbw_opamp_n_to_vbgtc:I left_hgbw_opamp_n_to_right_vref:I
*+ left_hgbw_opamp_n_to_vinref:I left_hgbw_opamp_n_to_gpio2_0[1:0]:I left_lp_opamp_p_to_gpio5_4[1:0]:I left_lp_opamp_p_to_dac0:I left_lp_opamp_p_to_analog0:I
*+ left_lp_opamp_p_to_amuxbusA:I right_instramp_p_to_left_rheostat2_out:I left_lp_opamp_p_to_sio0:I left_lp_opamp_p_to_left_vref:I left_lp_opamp_p_to_voutref:I
*+ left_lp_opamp_n_to_gpio5_5[1:0]:I left_lp_opamp_n_to_dac1:I left_lp_opamp_n_to_analog1:I left_lp_opamp_n_to_amuxbusB:I left_instramp_n_to_left_rheostat1_out:I
*+ left_lp_opamp_n_to_rheostat_tap:I left_lp_opamp_n_to_sio1:I left_lp_opamp_n_to_vbgsc:I left_lp_opamp_n_to_right_vref:I left_lp_opamp_n_to_vinref:I
*+ left_instramp_to_ulpcomp_p[1:0]:I left_instramp_to_comp_p[1:0]:I left_instramp_to_adc0[1:0]:I left_instramp_to_gpio4_4[1:0]:I left_instramp_to_analog1[1:0]:I
*+ left_instramp_to_amuxbusB[1:0]:I right_instramp_to_ulpcomp_n[1:0]:I right_instramp_to_comp_n[1:0]:I right_instramp_to_adc1[1:0]:I right_instramp_to_analog0[1:0]:I
*+ right_instramp_to_amuxbusA[1:0]:I right_instramp_to_gpio3_0[1:0]:I left_instramp_n_to_gpio5_7[1:0]:I left_instramp_n_to_analog1:I left_instramp_n_to_amuxbusB:I
*+ left_instramp_n_to_sio1:I left_instramp_n_to_right_vref:I left_instramp_n_to_vinref:I left_instramp_p_to_gpio5_6[1:0]:I left_instramp_p_to_analog0:I
*+ left_instramp_p_to_amuxbusA:I left_instramp_p_to_sio0:I left_instramp_p_to_tempsense:I left_instramp_p_to_left_vref:I left_instramp_p_to_voutref:I
*+ right_instramp_n_to_analog1:I right_instramp_n_to_amuxbusB:I right_instramp_n_to_sio1:I right_instramp_n_to_right_vref:I right_instramp_n_to_vinref:I
*+ right_instramp_n_to_gpio2_6[1:0]:I right_instramp_p_to_analog0:I right_instramp_p_to_amuxbusA:I right_instramp_p_to_tempsense:I right_instramp_p_to_left_vref:I
*+ right_instramp_p_to_voutref:I right_instramp_p_to_gpio2_7[1:0]:I ulpcomp_p_to_dac0:I ulpcomp_p_to_analog1:I ulpcomp_p_to_sio0:I ulpcomp_p_to_vbgtc:I
*+ ulpcomp_p_to_tempsense:I ulpcomp_p_to_left_vref:I ulpcomp_p_to_voutref:I ulpcomp_p_to_gpio6_0[1:0]:I ulpcomp_p_to_gpio1_7[1:0]:I ulpcomp_n_to_dac1:I
*+ ulpcomp_n_to_analog0:I ulpcomp_n_to_sio1:I ulpcomp_n_to_vbgsc:I ulpcomp_n_to_right_vref:I ulpcomp_n_to_vinref:I ulpcomp_n_to_gpio6_1[1:0]:I
*+ ulpcomp_n_to_gpio1_6[1:0]:I comp_p_to_dac0:I comp_p_to_analog1:I comp_p_to_sio0:I comp_p_to_vbgtc:I comp_p_to_tempsense:I comp_p_to_left_vref:I
*+ comp_p_to_voutref:I comp_p_to_gpio6_2[1:0]:I comp_p_to_gpio1_5[1:0]:I comp_n_to_dac1:I comp_n_to_analog0:I comp_n_to_sio1:I comp_n_to_vbgsc:I
*+ comp_n_to_right_vref:I comp_n_to_vinref:I comp_n_to_gpio6_3[1:0]:I comp_n_to_gpio1_4[1:0]:I adc0_to_dac0:I adc0_to_analog1:I adc0_to_vbgtc:I
*+ adc0_to_left_vref:I adc0_to_voutref:I adc0_to_gpio6_4[1:0]:I adc0_to_gpio1_3[1:0]:I adc1_to_dac1:I adc1_to_analog0:I adc1_to_vbgsc:I
*+ adc1_to_right_vref:I adc1_to_vinref:I adc1_to_gpio6_5[1:0]:I adc1_to_gpio1_2[1:0]:I sio0_connect[1:0]:I sio1_connect[1:0]:I analog0_connect[1:0]:I
*+ analog1_connect[1:0]:I vbgtc_to_user:I vbgsc_to_user:I user_to_comp_n[1:0]:I user_to_comp_p[1:0]:I user_to_ulpcomp_n[1:0]:I user_to_ulpcomp_p[1:0]:I
*+ user_to_adc0[1:0]:I user_to_adc1[1:0]:I dac0_to_user:I dac1_to_user:I tempsense_to_user:I right_vref_to_user:I left_vref_to_user:I vinref_to_user:I
*+ voutref_to_user:I adc0_to_tempsense:I user_adc0:I user_adc1:I user_comp_n:I user_comp_p:I user_ulpcomp_n:I user_ulpcomp_p:I user_voutref:O
*+ user_vinref:O user_left_vref:O user_right_vref:O user_tempsense:O user_dac0:O user_dac1:O user_vbgtc:O user_vbgsc:O user_gpio3_0_analog:B
*+ user_gpio3_1_analog:B user_gpio3_2_analog:B user_gpio3_3_analog:B user_gpio3_4_analog:B user_gpio3_5_analog:B user_gpio3_6_analog:B
*+ user_gpio3_7_analog:B user_gpio4_0_analog:B user_gpio4_1_analog:B user_gpio4_2_analog:B user_gpio4_3_analog:B user_gpio4_4_analog:B
*+ user_gpio4_5_analog:B user_gpio4_6_analog:B user_gpio4_7_analog:B gpio1_0:B gpio1_1:B gpio1_2:B gpio1_3:B gpio1_4:B gpio1_5:B gpio1_6:B gpio1_7:B
*+ gpio2_0:B gpio2_1:B gpio2_2:B gpio2_3:B gpio2_4:B gpio2_5:B gpio2_6:B gpio2_7:B gpio3_0:B gpio3_1:B gpio3_2:B gpio3_3:B gpio3_4:B gpio3_5:B
*+ gpio3_6:B gpio3_7:B gpio4_0:B gpio4_1:B gpio4_2:B gpio4_3:B gpio4_4:B gpio4_5:B gpio4_6:B gpio4_7:B gpio5_0:B gpio5_1:B gpio5_2:B gpio5_3:B
*+ gpio5_4:B gpio5_5:B gpio5_6:B gpio5_7:B gpio6_0:B gpio6_1:B gpio6_2:B gpio6_3:B gpio6_4:B gpio6_5:B gpio6_6:B gpio6_7:B analog0:B analog1:B
*+ sio0:B sio1:B voutref:I vinref:I right_vref:I left_vref:I vbg:O ibias_lsxo:O ibias_hsxo:O user_ibias50:O user_ibias100:O vccd0:B vssd0:B
*+ amuxbus_a_n:B amuxbus_b_n:B right_instramp_p_to_sio0:I dac0_to_analog1:I dac1_to_analog0:I audiodac_out_to_analog1[1:0]:I
*+ audiodac_outb_to_analog0[1:0]:I audiodac_inb:I bandgap_sel:I vddio:B vssio:B ldo_ref_sel:I tempsense_sel:I brownout_ena:I brownout_vtrip[2:0]:I
*+ brownout_otrip[2:0]:I brownout_isrc_sel:I brownout_oneshot:I brownout_rc_ena:I brownout_rc_dis:I brownout_vunder:O brownout_timeout:O brownout_filt:O
*+ brownout_unfilt:O
X1 vbgpwr vssio bandgap_trim[0] vcmosref net1 bandgap_trim[1] bandgap_trim[2] bandgap_trim[3] vccd0 vssd0 bandgap_ena vbgsc vbgtc
+ sky130_ak_ip__cmos_vref
x2 vccd0 vdda0 vssa0 comp_p comp_out comp_n comp_ena comp_hyst[1] comp_hyst[0] comp_trim[5] comp_trim[4] comp_trim[3] comp_trim[2]
+ comp_trim[1] comp_trim[0] ibias_comp vssd0 sky130_ak_ip__comparator
x3 vddio vbgpwr vssio ldo_ena vbg ldo_ref_sel vccd0 vssd0 sky130_am_ip__ldo_01v8
x9 adc1_dac_val[0] adc1_dac_val[1] adc1_dac_val[2] adc1_dac_val[3] adc1_dac_val[4] adc1_dac_val[5] adc1_dac_val[6] adc1_dac_val[7]
+ adc1_dac_val[8] adc1_dac_val[9] vdda0 vccd0 vssd0 vssa0 adc_vrefH adc_vrefL net27 adc1_reset net24 adc1_dac_val[10] adc1_dac_val[11] left_vref
+ vinref adc1 adc1_hold sky130_ef_ip__cdac3v_12bit
x10 vccd0 vssa0 vssd0 vdda0 left_rheostat1_b[0] left_rheostat1_in left_rheostat1_b[1] left_rheostat1_b[2] left_rheostat1_b[3]
+ left_rheostat1_tap left_rheostat1_b[4] left_rheostat1_b[5] left_rheostat1_b[6] left_rheostat1_b[7] left_hgbw_opamp_out sky130_ef_ip__rheostat_8bit
x12 vccd0 vdda0 ulpcomp_ena ulpcomp_out ulpcomp_n ulpcomp_p ulpcomp_clk vssd0 vssa0 sky130_icrg_ip__ulpcomp2
x14 net2 vccd0 vssd0 vbg tempsense_ena net3 sky130_od_ip__tempsensor_ext_vp
x17 overvoltage_out overvoltage_trim[0] vssd0 vssa0 vdda0 vccd0 ibias_ov vbg overvoltage_ena overvoltage_trim[3]
+ overvoltage_trim[2] overvoltage_trim[1] sky130_vbl_ip__overvoltage
x18 vssa1 vssa1 vssa1 vssa1 vssa1 vssa1 net9 net10 net11 net12 net13 net14 porb_h[0] net22 vccd0 vccd0 vdda1 vdda1_pwr_good
+ vccd1_pwr_good vccd1 vssa1 vssd0 vssd1 sky130_fd_io__top_pwrdetv2
x20 vccd0 vssa0 vssd0 vdda0 left_rheostat2_b[0] left_rheostat2_in left_rheostat2_b[1] left_rheostat2_b[2] left_rheostat2_b[3]
+ left_rheostat2_tap left_rheostat2_b[4] left_rheostat2_b[5] left_rheostat2_b[6] left_rheostat2_b[7] left_lp_opamp_out sky130_ef_ip__rheostat_8bit
x22 vccd0 vssa0 vssd0 vdda0 right_rheostat1_b[0] right_rheostat1_in right_rheostat1_b[1] right_rheostat1_b[2] right_rheostat1_b[3]
+ right_rheostat1_tap right_rheostat1_b[4] right_rheostat1_b[5] right_rheostat1_b[6] right_rheostat1_b[7] right_hgbw_opamp_out
+ sky130_ef_ip__rheostat_8bit
x24 vccd0 vssa0 vssd0 vdda0 right_rheostat2_b[0] right_rheostat2_in right_rheostat2_b[1] right_rheostat2_b[2] right_rheostat2_b[3]
+ right_rheostat2_tap right_rheostat2_b[4] right_rheostat2_b[5] right_rheostat2_b[6] right_rheostat2_b[7] right_lp_opamp_out
+ sky130_ef_ip__rheostat_8bit
x27 vssa2 vssa2 vssa2 vssa2 vssa2 vssa2 net15 net16 net17 net18 net19 net20 porb_h[0] net21 vccd0 vccd0 vdda2 vdda2_pwr_good
+ vccd2_pwr_good vccd2 vssa2 vssd0 vssd2 sky130_fd_io__top_pwrdetv2
x13 vccd0 vssa0 vssd0 vdda0 rdac1_value[0] dac_vrefH rdac1_value[1] rdac1_value[2] rdac1_value[3] dac1 rdac1_value[4]
+ rdac1_value[5] rdac1_ena rdac1_value[6] rdac1_value[7] dac_vrefL sky130_ef_ip__rdac3v_8bit
x29 vccd0 vssa0 vssd0 vdda0 rdac0_value[0] dac_vrefH rdac0_value[1] rdac0_value[2] rdac0_value[3] dac0 rdac0_value[4]
+ rdac0_value[5] rdac0_ena rdac0_value[6] rdac0_value[7] dac_vrefL sky130_ef_ip__rdac3v_8bit
x30 adc0_dac_val[0] adc0_dac_val[1] adc0_dac_val[2] adc0_dac_val[3] adc0_dac_val[4] adc0_dac_val[5] adc0_dac_val[6]
+ adc0_dac_val[7] adc0_dac_val[8] adc0_dac_val[9] vdda0 vccd0 vssd0 vssa0 adc_vrefH adc_vrefL net26 adc0_reset net23 adc0_dac_val[10]
+ adc0_dac_val[11] right_vref voutref adc0 adc0_hold sky130_ef_ip__cdac3v_12bit
x33 vdda0 vccd0 vssd0 vssa0 adc1 comp_n ulpcomp_n right_instramp_to_ulpcomp_n[1] right_instramp_to_ulpcomp_n[0] right_instramp_out
+ right_hgbw_opamp_to_ulpcomp_n[1] right_hgbw_opamp_to_ulpcomp_n[0] right_lp_opamp_to_ulpcomp_p[1] right_lp_opamp_to_ulpcomp_p[0] left_lp_opamp_to_ulpcomp_n[1]
+ left_lp_opamp_to_ulpcomp_n[0] left_hgbw_opamp_to_ulpcomp_p[1] left_hgbw_opamp_to_ulpcomp_p[0] left_instramp_to_ulpcomp_p[1] left_instramp_to_ulpcomp_p[0]
+ right_hgbw_opamp_out right_instramp_to_comp_n[1] right_instramp_to_comp_n[0] right_hgbw_opamp_to_comp_n[1] right_hgbw_opamp_to_comp_n[0]
+ right_lp_opamp_to_comp_p[1] right_lp_opamp_to_comp_p[0] left_lp_opamp_to_comp_n[1] left_lp_opamp_to_comp_n[0] left_hgbw_opamp_to_comp_p[1]
+ left_hgbw_opamp_to_comp_p[0] left_instramp_to_comp_p[1] left_instramp_to_comp_p[0] right_lp_opamp_out right_instramp_to_adc1[1] right_instramp_to_adc1[0]
+ right_hgbw_opamp_to_adc1[1] right_hgbw_opamp_to_adc1[0] right_lp_opamp_to_adc0[1] right_lp_opamp_to_adc0[0] left_lp_opamp_to_adc1[1] left_lp_opamp_to_adc1[0]
+ left_hgbw_opamp_to_adc0[1] left_hgbw_opamp_to_adc0[0] left_lp_opamp_out left_instramp_to_adc0[1] left_instramp_to_adc0[0] left_hgbw_opamp_out
+ left_instramp_out adc0 ulpcomp_p comp_p switch_array_18
x34 vdda0 vccd0 vssd0 vssa0 right_instramp_to_amuxbusA[1] right_instramp_to_amuxbusA[0] right_instramp_out
+ left_hgbw_opamp_to_amuxbusB[1] left_hgbw_opamp_to_amuxbusB[0] left_lp_opamp_to_amuxbusA[1] left_lp_opamp_to_amuxbusA[0] right_lp_opamp_to_amuxbusB[1]
+ right_lp_opamp_to_amuxbusB[0] right_hgbw_opamp_to_amuxbusA[1] right_hgbw_opamp_to_amuxbusA[0] left_instramp_to_amuxbusB[1] left_instramp_to_amuxbusB[0]
+ right_hgbw_opamp_out right_instramp_to_analog0[1] right_instramp_to_analog0[0] left_hgbw_opamp_to_analog1[1] left_hgbw_opamp_to_analog1[0]
+ left_lp_opamp_to_analog0[1] left_lp_opamp_to_analog0[0] right_lp_opamp_to_analog1[1] right_lp_opamp_to_analog1[0] right_hgbw_opamp_to_analog0[1]
+ right_hgbw_opamp_to_analog0[0] left_instramp_to_analog1[1] left_instramp_to_analog1[0] right_lp_opamp_out left_lp_opamp_out left_hgbw_opamp_out
+ left_instramp_out analog1 analog1_core analog0 analog0_core amuxbus_b_n amuxbus_a_n analog1_connect[1] analog1_connect[0] analog0_connect[1]
+ analog0_connect[0] switch_array_14
x35 vdda0 vccd0 vssd0 vssa0 gpio4_4 left_instramp_to_gpio4_4[1] left_instramp_to_gpio4_4[0] left_instramp_out
+ left_hgbw_opamp_to_gpio4_5[1] left_hgbw_opamp_to_gpio4_5[0] right_lp_opamp_to_gpio4_7[1] right_lp_opamp_to_gpio4_7[0] right_hgbw_opamp_to_gpio4_6[1]
+ right_hgbw_opamp_to_gpio4_6[0] gpio4_5 left_hgbw_opamp_out gpio4_7 right_lp_opamp_out gpio4_6 right_hgbw_opamp_out switch_array_4
x36 vdda0 vccd0 vssd0 vssa0 gpio4_0 left_lp_opamp_to_gpio4_0[1] left_lp_opamp_to_gpio4_0[0] left_lp_opamp_out
+ left_hgbw_opamp_to_gpio4_1[1] left_hgbw_opamp_to_gpio4_1[0] right_lp_opamp_to_gpio4_3[1] right_lp_opamp_to_gpio4_3[0] right_hgbw_opamp_to_gpio4_2[1]
+ right_hgbw_opamp_to_gpio4_2[0] gpio4_1 left_hgbw_opamp_out gpio4_3 right_lp_opamp_out gpio4_2 right_hgbw_opamp_out switch_array_4
x37 vdda0 vccd0 vssd0 vssa0 gpio3_4 left_lp_opamp_to_gpio3_4[1] left_lp_opamp_to_gpio3_4[0] left_lp_opamp_out
+ left_hgbw_opamp_to_gpio3_5[1] left_hgbw_opamp_to_gpio3_5[0] right_lp_opamp_to_gpio3_7[1] right_lp_opamp_to_gpio3_7[0] right_hgbw_opamp_to_gpio3_6[1]
+ right_hgbw_opamp_to_gpio3_6[0] gpio3_5 left_hgbw_opamp_out gpio3_7 right_lp_opamp_out gpio3_6 right_hgbw_opamp_out switch_array_4
x38 vdda0 vccd0 vssd0 vssa0 gpio3_3 right_lp_opamp_to_gpio3_3[1] right_lp_opamp_to_gpio3_3[0] right_lp_opamp_out
+ right_hgbw_opamp_to_gpio3_2[1] right_hgbw_opamp_to_gpio3_2[0] right_instramp_to_gpio3_0[1] right_instramp_to_gpio3_0[0] left_hgbw_opamp_to_gpio3_1[1]
+ left_hgbw_opamp_to_gpio3_1[0] gpio3_2 right_hgbw_opamp_out gpio3_0 right_instramp_out gpio3_1 left_hgbw_opamp_out switch_array_4
x39 vdda0 vccd0 vssd0 vssa0 gpio5_5 left_lp_opamp_n_to_gpio5_5[1] left_lp_opamp_n_to_gpio5_5[0] left_lp_opamp_in_n
+ left_lp_opamp_p_to_gpio5_4[1] left_lp_opamp_p_to_gpio5_4[0] left_instramp_p_to_gpio5_6[1] left_instramp_p_to_gpio5_6[0] left_instramp_n_to_gpio5_7[1]
+ left_instramp_n_to_gpio5_7[0] gpio5_4 left_lp_opamp_in_p gpio5_6 left_instramp_in_p gpio5_7 left_instramp_in_n switch_array_4
x40 vdda0 vccd0 vssd0 vssa0 gpio6_1 ulpcomp_n_to_gpio6_1[1] ulpcomp_n_to_gpio6_1[0] ulpcomp_n ulpcomp_p_to_gpio6_0[1]
+ ulpcomp_p_to_gpio6_0[0] comp_p_to_gpio6_2[1] comp_p_to_gpio6_2[0] comp_n_to_gpio6_3[1] comp_n_to_gpio6_3[0] gpio6_0 ulpcomp_p gpio6_2 comp_p gpio6_3
+ comp_n switch_array_4
x41 vdda0 vccd0 vssd0 vssa0 gpio6_5 adc1_to_gpio6_5[1] adc1_to_gpio6_5[0] adc1 adc0_to_gpio6_4[1] adc0_to_gpio6_4[0]
+ adc_refh_to_gpio6_6[1] adc_refh_to_gpio6_6[0] adc_refl_to_gpio6_7[1] adc_refl_to_gpio6_7[0] gpio6_4 adc0 gpio6_6 adc_vrefH gpio6_7 adc_vrefL
+ switch_array_4
x42 vdda0 vccd0 vssd0 vssa0 gpio5_1 right_hgbw_opamp_n_to_gpio5_1[1] right_hgbw_opamp_n_to_gpio5_1[0] right_hgbw_opamp_in_n
+ right_hgbw_opamp_p_to_gpio5_0[1] right_hgbw_opamp_p_to_gpio5_0[0] left_hgbw_opamp_p_to_gpio5_2[1] left_hgbw_opamp_p_to_gpio5_2[0] left_hgbw_opamp_n_to_gpio5_3[1]
+ left_hgbw_opamp_n_to_gpio5_3[0] gpio5_0 right_hgbw_opamp_in_p gpio5_2 left_hgbw_opamp_in_p gpio5_3 left_hgbw_opamp_in_n switch_array_4
x43 vdda0 vccd0 vssd0 vssa0 gpio2_2 right_hgbw_opamp_n_to_gpio2_2[1] right_hgbw_opamp_n_to_gpio2_2[0] right_hgbw_opamp_in_n
+ right_hgbw_opamp_p_to_gpio2_3[1] right_hgbw_opamp_p_to_gpio2_3[0] dac_refl_to_gpio1_0[1] dac_refl_to_gpio1_0[0] dac_refh_to_gpio1_1[1] dac_refh_to_gpio1_1[0]
+ gpio2_3 right_hgbw_opamp_in_p gpio1_0 dac_vrefL gpio1_1 dac_vrefH switch_array_4
x44 vdda0 vccd0 vssd0 vssa0 gpio1_6 ulpcomp_n_to_gpio1_6[1] ulpcomp_n_to_gpio1_6[0] ulpcomp_n ulpcomp_p_to_gpio1_7[1]
+ ulpcomp_p_to_gpio1_7[0] left_hgbw_opamp_n_to_gpio2_0[1] left_hgbw_opamp_n_to_gpio2_0[0] left_hgbw_opamp_p_to_gpio2_1[1] left_hgbw_opamp_p_to_gpio2_1[0]
+ gpio1_7 ulpcomp_p gpio2_0 left_hgbw_opamp_in_n gpio2_1 left_hgbw_opamp_in_p switch_array_4
x45 vdda0 vccd0 vssd0 vssa0 gpio1_2 adc1_to_gpio1_2[1] adc1_to_gpio1_2[0] adc1 adc0_to_gpio1_3[1] adc0_to_gpio1_3[0]
+ comp_n_to_gpio1_4[1] comp_n_to_gpio1_4[0] comp_p_to_gpio1_5[1] comp_p_to_gpio1_5[0] gpio1_3 adc0 gpio1_4 comp_n gpio1_5 comp_p switch_array_4
x46 vdda0 vccd0 vssd0 vssa0 gpio2_7 right_instramp_p_to_gpio2_7[1] right_instramp_p_to_gpio2_7[0] right_instramp_in_p
+ right_instramp_n_to_gpio2_6[1] right_instramp_n_to_gpio2_6[0] right_lp_opamp_p_to_gpio2_5[1] right_lp_opamp_p_to_gpio2_5[0] right_lp_opamp_n_to_gpio2_4[1]
+ right_lp_opamp_n_to_gpio2_4[0] gpio2_6 right_instramp_in_n gpio2_5 right_lp_opamp_in_p gpio2_4 right_lp_opamp_in_n switch_array_4
* noconn rdac0_value[11:8]
* noconn rdac1_value[11:8]
* noconn adc0_dac_val[15:12]
* noconn adc1_dac_val[15:12]
x47 vdda0 vssa0 vccd0 vssd0 analog1_core amuxbus_a_n amuxbus_b_n analog0_core right_instramp_n_to_analog1
+ right_instramp_p_to_amuxbusA right_instramp_n_to_amuxbusB right_instramp_p_to_analog0 right_instramp_in_n right_hgbw_opamp_n_to_analog1 right_instramp_in_p
+ right_hgbw_opamp_n_to_amuxbusB right_hgbw_opamp_p_to_amuxbusA right_hgbw_opamp_p_to_analog0 right_hgbw_opamp_in_n right_hgbw_opamp_in_p right_lp_opamp_in_n
+ right_lp_opamp_in_p right_lp_opamp_n_to_analog1 right_lp_opamp_p_to_amuxbusA right_lp_opamp_p_to_analog0 right_lp_opamp_n_to_amuxbusB
+ left_instramp_in_n left_instramp_in_p left_hgbw_opamp_in_n left_hgbw_opamp_in_p left_lp_opamp_n_to_analog1 left_lp_opamp_p_to_amuxbusA
+ left_lp_opamp_n_to_amuxbusB left_lp_opamp_p_to_analog0 left_lp_opamp_in_n left_lp_opamp_in_p ulpcomp_p ulpcomp_n left_hgbw_opamp_n_to_analog1
+ left_hgbw_opamp_p_to_analog0 left_hgbw_opamp_n_to_amuxbusB left_hgbw_opamp_p_to_amuxbusA comp_p comp_n adc0 adc1 left_instramp_n_to_analog1 dac0
+ left_instramp_p_to_analog0 left_instramp_n_to_amuxbusB left_instramp_p_to_amuxbusA dac1 ulpcomp_p_to_analog1 ulpcomp_n_to_analog0 comp_p_to_analog1
+ comp_n_to_analog0 adc0_to_analog1 adc1_to_analog0 dac0_to_analog1 dac1_to_analog0 simple_switch_array_32
x48 vdda0 vssa0 vccd0 vssd0 vbgtc vbgsc left_vref tempsense_out right_vref voutref vinref right_instramp_p_to_left_vref
+ right_instramp_n_to_right_vref right_instramp_p_to_tempsense right_instramp_n_to_vinref right_instramp_p_to_voutref right_instramp_in_n right_instramp_in_p
+ right_hgbw_opamp_n_to_vbgsc right_hgbw_opamp_in_n right_hgbw_opamp_in_p right_hgbw_opamp_n_to_right_vref right_hgbw_opamp_p_to_left_vref
+ right_hgbw_opamp_n_to_vinref right_hgbw_opamp_p_to_voutref right_lp_opamp_in_n right_lp_opamp_in_p right_lp_opamp_n_to_vbgtc left_instramp_in_n
+ left_instramp_in_p right_lp_opamp_n_to_right_vref right_lp_opamp_p_to_left_vref right_lp_opamp_p_to_voutref right_lp_opamp_n_to_vinref
+ left_hgbw_opamp_in_n left_lp_opamp_n_to_vbgsc left_hgbw_opamp_in_p left_lp_opamp_in_n left_lp_opamp_in_p right_lp_opamp_p_to_tempsense
+ left_lp_opamp_n_to_right_vref left_lp_opamp_p_to_left_vref left_lp_opamp_p_to_voutref left_lp_opamp_n_to_vinref ulpcomp_p ulpcomp_n
+ left_hgbw_opamp_p_to_tempsense comp_p comp_n left_hgbw_opamp_n_to_right_vref left_hgbw_opamp_p_to_left_vref left_hgbw_opamp_p_to_voutref
+ left_hgbw_opamp_n_to_vinref adc0 adc1 left_instramp_n_to_right_vref left_instramp_p_to_tempsense left_instramp_p_to_left_vref left_instramp_p_to_voutref
+ left_instramp_n_to_vinref ulpcomp_p_to_vbgtc ulpcomp_n_to_vbgsc ulpcomp_n_to_vinref ulpcomp_p_to_left_vref ulpcomp_n_to_right_vref ulpcomp_p_to_tempsense
+ ulpcomp_p_to_voutref comp_p_to_vbgtc comp_n_to_vbgsc comp_n_to_vinref comp_p_to_left_vref comp_n_to_right_vref comp_p_to_tempsense comp_p_to_voutref
+ adc0_to_vbgtc adc1_to_vbgsc adc1_to_vinref adc1_to_right_vref adc0_to_left_vref adc0_to_tempsense adc0_to_voutref left_hgbw_opamp_n_to_vbgtc
+ simple_switch_array_53
x49 vdda0 vssa0 vccd0 vssd0 right_hgbw_opamp_n_to_dac1 right_hgbw_opamp_p_to_dac0 right_hgbw_opamp_in_n right_hgbw_opamp_in_p
+ right_lp_opamp_n_to_dac1 right_lp_opamp_p_to_dac0 right_lp_opamp_in_n right_lp_opamp_in_p left_hgbw_opamp_in_n left_hgbw_opamp_in_p
+ left_lp_opamp_n_to_dac1 left_lp_opamp_p_to_dac0 left_lp_opamp_in_n left_lp_opamp_in_p ulpcomp_p ulpcomp_n left_hgbw_opamp_n_to_dac1
+ left_hgbw_opamp_p_to_dac0 comp_p comp_n adc0 adc1 ulpcomp_n_to_dac1 ulpcomp_p_to_dac0 dac0 dac1 comp_n_to_dac1 comp_p_to_dac0 adc1_to_dac1 adc0_to_dac0
+ simple_switch_array_14
x50 vdda0 vssa0 vccd0 vssd0 right_instramp_n_to_sio1 right_instramp_p_to_sio0 sio0_core sio1_core right_hgbw_opamp_n_to_sio1
+ right_hgbw_opamp_p_to_sio0 right_instramp_in_n right_instramp_in_p right_hgbw_opamp_in_n right_hgbw_opamp_in_p right_lp_opamp_n_to_sio1 right_lp_opamp_in_n
+ right_lp_opamp_p_to_sio0 right_lp_opamp_in_p left_instramp_in_n left_instramp_in_p left_hgbw_opamp_in_n left_lp_opamp_n_to_sio1 left_lp_opamp_p_to_sio0
+ left_hgbw_opamp_in_p left_lp_opamp_in_n left_lp_opamp_in_p ulpcomp_p left_hgbw_opamp_n_to_sio1 left_hgbw_opamp_p_to_sio0 ulpcomp_n comp_p comp_n
+ left_instramp_n_to_sio1 left_instramp_p_to_sio0 ulpcomp_n_to_sio1 ulpcomp_p_to_sio0 comp_n_to_sio1 comp_p_to_sio0 simple_switch_array_16
x51 user_to_comp_n[1] user_to_comp_n[0] user_to_comp_p[1] user_to_comp_p[0] vdda0 user_to_ulpcomp_n[1] user_to_ulpcomp_n[0] vssa0
+ vccd0 user_to_ulpcomp_p[1] user_to_ulpcomp_p[0] vssd0 user_to_adc0[1] user_to_adc0[0] user_to_adc1[1] user_to_adc1[0] vbgtc_to_user
+ user_comp_n comp_n user_vbgtc vbgtc vbgsc_to_user user_comp_p comp_p user_vbgsc vbgsc dac0_to_user user_ulpcomp_n ulpcomp_n user_dac0 dac0
+ dac1_to_user user_ulpcomp_p ulpcomp_p user_dac1 dac1 tempsense_to_user user_adc0 adc0 user_tempsense tempsense_out right_vref_to_user
+ user_adc1 adc1 user_right_vref right_vref left_vref_to_user user_left_vref left_vref vinref_to_user user_vinref vinref voutref_to_user
+ user_voutref voutref user_switch_array_15
x52 vdda0 vssa0 vccd0 vssd0 right_instramp_p_to_right_rheostat1_out right_instramp_n_to_right_rheostat1_out right_rheostat1_in
+ right_hgbw_opamp_in_n left_instramp_p_to_left_rheostat1_out right_hgbw_opamp_n_to_rheostat_tap right_lp_opamp_in_n right_rheostat1_tap
+ left_hgbw_opamp_in_n right_instramp_p_to_left_rheostat2_out left_instramp_n_to_left_rheostat1_out left_lp_opamp_in_n right_rheostat2_in
+ right_lp_opamp_n_to_rheostat_tap left_instramp_p_to_right_rheostat2_out right_rheostat2_tap right_instramp_n_to_left_rheostat2_out left_rheostat2_in
+ left_lp_opamp_n_to_rheostat_tap left_rheostat2_tap left_instramp_n_to_right_rheostat2_out left_rheostat1_in left_hgbw_opamp_n_to_rheostat_tap left_rheostat1_tap
+ left_instramp_in_n left_instramp_in_p right_instramp_in_n right_instramp_in_p simple_switch_array_12
x53 vdda0 vccd0 vssd0 vssa0 gpio1_2 ibias_test_to_gpio1_2[1] ibias_test_to_gpio1_2[0] ibias_test vbg_test_to_gpio1_1[1]
+ vbg_test_to_gpio1_1[0] gpio1_1 vbg switch_array_2
x54 vdda0 vccd0 vssd0 vssa0 gpio1_3 idac_to_gpio1_3[1] idac_to_gpio1_3[0] idac_snk idac_to_gpio1_2[1] idac_to_gpio1_2[0] gpio1_2
+ idac_src switch_array_2
x55 vdda0 vccd0 vssd0 vssa0 sio1 sio1_connect[1] sio1_connect[0] sio1_core sio0_connect[1] sio0_connect[0] sio0 sio0_core
+ switch_array_2
x56 vdda0 vccd0 vssd0 vssa0 analog1_core audiodac_out_to_analog1[1] audiodac_out_to_analog1[0] audiodac_out
+ audiodac_outb_to_analog0[1] audiodac_outb_to_analog0[0] analog0_core audiodac_outb switch_array_2
x5 vssa0 tempsense_sel net2 vdda0 net3 tempsense_out vccd0 vssd0 simple_analog_mux_sel1v8
x6 vssa0 bandgap_sel net25 vdda0 vcmosref vbg vccd0 vssd0 simple_analog_mux_sel1v8
x7 idac_ena vdda1 vbg ibias_ref_select vccd0 vssd0 vdda0 idac_value[7] idac_value[6] idac_value[5] idac_value[4] idac_value[3]
+ idac_value[2] idac_value[1] idac_value[0] vssa0 idac_src idac_snk sky130_ef_ip__idac3v_8bit
* noconn idac_value[11:8]
x59 vdda0 vssa0 net8 vccd0 net7 vssd0 brownout_unfilt vbg brownout_otrip[2] brownout_otrip[1] brownout_otrip[0] net6 brownout_filt
+ brownout_vtrip[2] brownout_vtrip[1] brownout_vtrip[0] net5 brownout_ena brownout_rc_ena net4 brownout_rc_dis brownout_timeout brownout_vunder
+ brownout_oneshot brownout_isrc_sel brownout_ibias sky130_ajc_ip__brownout
* noconn #net7
* noconn #net8
* noconn #net6
* noconn #net5
* noconn #net4
* noconn #net9
* noconn #net10
* noconn #net11
* noconn #net12
* noconn #net13
* noconn #net14
* noconn #net15
* noconn #net16
* noconn #net17
* noconn #net18
* noconn #net19
* noconn #net20
* noconn #net22
* noconn #net21
* noconn ibias_idac
* noconn #net1
R15 gpio3_0 user_gpio3_0_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R1 gpio3_1 user_gpio3_1_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R2 gpio3_2 user_gpio3_2_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R3 gpio3_3 user_gpio3_3_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R4 gpio3_4 user_gpio3_4_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R5 gpio3_5 user_gpio3_5_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R6 gpio3_6 user_gpio3_6_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R7 gpio3_7 user_gpio3_7_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R8 gpio4_0 user_gpio4_0_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R9 gpio4_1 user_gpio4_1_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R10 gpio4_2 user_gpio4_2_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R11 gpio4_3 user_gpio4_3_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R12 gpio4_4 user_gpio4_4_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R13 gpio4_5 user_gpio4_5_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R14 gpio4_6 user_gpio4_6_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
R16 gpio4_7 user_gpio4_7_analog sky130_fd_pr__res_generic_m4 W=1 L=1 m=1
XC1 vbgpwr vssio sky130_fd_pr__cap_mim_m3_2 W=10 L=10 m=18
XC2 vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 m=35
XC3 vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 m=20
XC4 vccd0 vssd0 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 m=10
XC5 vddio vssio sky130_fd_pr__cap_mim_m3_2 W=10 L=10 m=32
x26 audiodac_out vdda0 vccd0 audiodac_in audiodac_inb vssa0 audiodac_outb sky130_iic_ip__audiodac_drv_lite
XC6 vcmosref vssio sky130_fd_pr__cap_mim_m3_2 W=10 L=10 m=10
* noconn #net23
* noconn #net24
x28 left_instramp_G2[4] left_instramp_G2[3] left_instramp_G2[2] left_instramp_G2[1] left_instramp_G2[0] left_instramp_G1[4]
+ left_instramp_G1[3] left_instramp_G1[2] left_instramp_G1[1] left_instramp_G1[0] left_vref ibias_instr1 vdda0 left_instramp_in_n vccd0
+ left_instramp_out vssa0 vssd0 left_instramp_in_p sky130_pa_ip__instramp
x58 right_instramp_G2[4] right_instramp_G2[3] right_instramp_G2[2] right_instramp_G2[1] right_instramp_G2[0] right_instramp_G1[4]
+ right_instramp_G1[3] right_instramp_G1[2] right_instramp_G1[1] right_instramp_G1[0] right_vref ibias_instr2 vdda0 right_instramp_in_n vccd0
+ right_instramp_out vssa0 vssd0 right_instramp_in_p sky130_pa_ip__instramp
* noconn right_instramp_ena
* noconn left_instramp_ena
x19 adc1_comp_out vccd0 vssd0 vdda0 vssa0 net27 left_vref adc1_ena sky130_ef_ip__scomp3v
x8 adc0_comp_out vccd0 vssd0 vdda0 vssa0 net26 right_vref adc0_ena sky130_ef_ip__scomp3v
x11 vdda0 left_hgbw_opamp_out left_hgbw_opamp_ibias left_hgbw_opamp_in_n left_hgbw_opamp_in_p vssa0 vccd0 vssd0
+ left_hgbw_opamp_ena sky130_td_ip__opamp_hp_narrow
x31 vdda0 left_lp_opamp_out left_lp_opamp_ibias left_lp_opamp_in_n left_lp_opamp_in_p vssa0 vccd0 vssd0 left_lp_opamp_ena
+ sky130_td_ip__opamp_hp_narrow
x32 vdda0 right_lp_opamp_out right_lp_opamp_ibias right_lp_opamp_in_n right_lp_opamp_in_p vssa0 vccd0 vssd0 right_lp_opamp_ena
+ sky130_td_ip__opamp_hp_narrow
x60 vdda0 right_hgbw_opamp_out right_hgbw_opamp_ibias right_hgbw_opamp_in_n right_hgbw_opamp_in_p vssa0 vccd0 vssd0
+ right_hgbw_opamp_ena sky130_td_ip__opamp_hp_narrow
x16 vccd0 net25 vssd0 bandgap_ibias bandgap_trim[15] bandgap_trim[14] bandgap_trim[13] bandgap_trim[12] bandgap_trim[11]
+ bandgap_trim[10] bandgap_trim[9] bandgap_trim[8] bandgap_trim[7] bandgap_trim[6] bandgap_trim[5] bandgap_trim[4] bandgap_trim[3] bandgap_trim[2]
+ bandgap_trim[1] bandgap_trim[0] vssd0 sky130_cw_ip__bandgap_nobias
x4 ibias_ena vdda0 vssa0 vdda1 vccd0 vbg ibias_ref_select vssd0 left_lp_opamp_ibias ibias_src_ena[0] ibias_src_ena[1]
+ ibias_src_ena[2] right_lp_opamp_ibias ibias_src_ena[3] ibias_src_ena[4] left_hgbw_opamp_ibias ibias_src_ena[5] right_hgbw_opamp_ibias
+ ibias_src_ena[6] ibias_src_ena[7] ibias_instr1 ibias_src_ena[8] ibias_src_ena[9] ibias_instr2 ibias_src_ena[10] ibias_src_ena[11] ibias_lsxo
+ ibias_src_ena[12] ibias_hsxo ibias_src_ena[13] ibias_src_ena[14] ibias_snk_ena[0] ibias_comp ibias_src_ena[15] ibias_src_ena[16] ibias_snk_ena[1]
+ ibias_ov ibias_src_ena[17] ibias_src_ena[18] ibias_idac ibias_src_ena[19] brownout_ibias ibias_src_ena[20] user_ibias50 ibias_src_ena[21]
+ user_ibias100 ibias_src_ena[22] ibias_snk_ena[2] ibias_src_ena[23] ibias_test ibias_snk_ena[3] bandgap_ibias sky130_ef_ip__biasgen4
x21 por vssio vddio vccd0 porb vssd0 porb_h[1] porb_h[0] sky130_sw_ip__por
.ends

* expanding   symbol:  sky130_ak_ip__cmos_vref.sym # of pins=13
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ak_ip__cmos_vref/xschem/sky130_ak_ip__cmos_vref.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ak_ip__cmos_vref/xschem/sky130_ak_ip__cmos_vref.sch
.subckt sky130_ak_ip__cmos_vref avdd18 avss trim0 vbg vptat trim1 trim2 trim3 dvdd dvss ena vbgsc vbgtg
*.PININFO vbg:O avss:B avdd18:B dvss:B ena:I vbgsc:O vbgtg:O trim3:I trim2:I trim1:I trim0:I vptat:O dvdd:B
XM2 vref vref vptat avss sky130_fd_pr__nfet_01v8 L=10 W=2 nf=1 m=1
XM1 vptat vref avss avss sky130_fd_pr__nfet_01v8 L=20 W=2.5 nf=1 m=1
XM9 vref pbias net5 avdd_ena sky130_fd_pr__pfet_01v8 L=10 W=50 nf=4 m=1
XM20 avdd_ena net11 avdd18 dvdd sky130_fd_pr__pfet_01v8 L=0.3 W=10 nf=1 m=1
x1 net4 pbias vref vptat avss sbvfcm
x2 avdd_ena vbg vref net1 net2 avss output_amp
XM3 net2 pbias net3 avdd_ena sky130_fd_pr__pfet_01v8 L=10 W=5 nf=1 m=1
Vm_b1 avdd_ena net5 0
.save i(vm_b1)
Vm_b2 avdd_ena net4 0
.save i(vm_b2)
Vm_b3 avdd_ena net3 0
.save i(vm_b3)
x3 net6 net10 net8 net7 net9 avss trim_res
XR4 net6 net1 avss sky130_fd_pr__res_xhigh_po_0p69 L=264.5 mult=1 m=1
XR3 net1 vbgsc avss sky130_fd_pr__res_xhigh_po_0p69 L=74.5 mult=1 m=1
XR2 vbgsc vbgtg avss sky130_fd_pr__res_xhigh_po_0p69 L=8.6 mult=1 m=1
XR1 vbgtg vbg avss sky130_fd_pr__res_xhigh_po_0p69 L=54.5 mult=1 m=1
x5 trim3 dvss dvss dvdd dvdd net7 sky130_fd_sc_hd__buf_1
x6 trim2 dvss dvss dvdd dvdd net8 sky130_fd_sc_hd__buf_1
x7 trim1 dvss dvss dvdd dvdd net9 sky130_fd_sc_hd__buf_1
x8 trim0 dvss dvss dvdd dvdd net10 sky130_fd_sc_hd__buf_1
x9 trim0 dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
x14 ena dvss dvss dvdd dvdd net11 sky130_fd_sc_hd__inv_2
x4 trim1 dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
x10 trim2 dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
x11 trim3 dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
x12 ena dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
x13 dvss dvss dvdd dvdd sky130_fd_sc_hd__decap_6
.ends


* expanding   symbol:  sky130_ak_ip__comparator.sym # of pins=11
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ak_ip__comparator/xschem/sky130_ak_ip__comparator.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ak_ip__comparator/xschem/sky130_ak_ip__comparator.sch
.subckt sky130_ak_ip__comparator DVDD AVDD AGND Vinp Vout Vinm en hyst[1] hyst[0] trim[5] trim[4] trim[3] trim[2] trim[1] trim[0]
+ ibias DGND
*.PININFO Vinp:I Vinm:I AVDD:I AGND:I en:I hyst[1:0]:I trim[5:0]:I Vout:O DGND:I ibias:I DVDD:I
XM7 bias_n bias_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=2
XM6 Vfold_p Vinm Vxm AGND sky130_fd_pr__nfet_g5v0d10v5 L=1.5 W=8 nf=1 m=28
XM2 net1 bias_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=48
XM1 Vfold_m Vinp Vxm AGND sky130_fd_pr__nfet_g5v0d10v5 L=1.5 W=8 nf=1 m=28
XM4 net4 bias_var_tailp AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=96
XM5 Vfold_bot_p Vinm Vxp AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1.5 W=8 nf=1 m=28
XM17 Vfold_bot_m Vinp Vxp AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1.5 W=8 nf=1 m=28
XM22 net2 bias_stg2 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=4
XM23 Vom_stg2 Vop net2 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM24 Vop_stg2 Vom net2 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM25 Vop_stg2 Vop_stg2 AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM26 Vom_stg2 Vom_stg2 AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM27 net3 Vom_stg2 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM28 Vdiff Vop_stg2 DGND DGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM29 Vdiff net3 DVDD DVDD sky130_fd_pr__pfet_01v8 L=1 W=4 nf=1 m=2
XM30 net3 net3 DVDD DVDD sky130_fd_pr__pfet_01v8 L=1 W=4 nf=1 m=2
XM31 Vout_int Vdiff DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM44 Vout_int Vdiff DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM45 net52 ibias bias_n AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=1
XM48 bias_n enb_hv AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=4
XM40 net11 bias_n net5 AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=8
XM53 Vfold_p Voutb Vx_hyst_n AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=8
XM54 Vfold_m Vout_int Vx_hyst_n AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=8
XM73 net12 bias_n net24 AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=3
XM75 Voutb Vout_int DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM76 Voutb Vout_int DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM90 Vxm casc_n net1 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=48
XM91 Vxp casc_p net4 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=96
XM94 net10 bias_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=2
XM95 bias_p bias_p AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=4
XM16 net5 hyst1_hv AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=8
XM33 net24 hyst0_hv AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=3
XM67 Vop_stg2 Vom_stg2 AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=2 W=0.5 nf=1 m=1
XM69 Vom_stg2 Vop_stg2 AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=2 W=0.5 nf=1 m=1
XM15 bias_p en_hv AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=2 m=4
x2 AVDD trim2b_hv trim2_hv trim[2] AGND DVDD DGND level_shifter_up
x4 AVDD trim1b_hv trim1_hv trim[1] AGND DVDD DGND level_shifter_up
x5 AVDD trim0b_hv trim0_hv trim[0] AGND DVDD DGND level_shifter_up
x6 AVDD enb_hv en_hv en AGND DVDD DGND level_shifter_up
x7 AVDD hyst1b_hv hyst1_hv hyst[1] AGND DVDD DGND level_shifter_up
x8 AVDD hyst0b_hv hyst0_hv hyst[0] AGND DVDD DGND level_shifter_up
XM32 Vdiff enb_hv DGND DGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=4
XM34 casc_n bias_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=2
XM36 AVDD ibias casc_n AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM3 Vfold_bot_p Vom AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=12
XM9 Vfold_p bias_p AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=24
XM10 Vfold_p bias_var_p AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=56
XM13 Vfold_bot_p bias_var_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=28
XM19 Vop casc_p Vfold_p AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=80
XM21 Vop casc_n Vfold_bot_p AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=40
XM38 net7 Vinm net6 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1.5 W=8 nf=1 m=1
XM39 net7 Vinp net6 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1.5 W=8 nf=1 m=1
XM49 net7 bias_var_p AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=4
XM60 net9 bias_var_p AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=4
XM61 net8 bias_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=2
XM62 net50 bias_var_tailp AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=4
XM68 net48 bias_var_tailp AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=4
XM70 bias_var_n bias_var_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=2
XM8 Vfold_bot_m bias_var_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=28
XM11 Vfold_m bias_var_p AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=56
XM12 Vfold_m bias_p AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=24
XM14 Vfold_bot_m Vom AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=12
XM18 Vom casc_p Vfold_m AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=80
XM20 Vom casc_n Vfold_bot_m AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=40
XM84 bias_var_tailp casc_n net8 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM85 bias_var_tailp casc_p net9 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM86 bias_p casc_n net10 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM88 Vx_hyst_n casc_n net11 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=8
XM89 Vfold_m net35 net29 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1.5 W=8 nf=1 m=4
XM92 net13 bias_var_tailn AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=6
XM93 Vfold_p net34 net29 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1.5 W=8 nf=1 m=4
XM97 net29 casc_n net13 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=6
x1 AVDD trim3b_hv trim3_hv trim[3] AGND DVDD DGND level_shifter_up
XM63 net21 bias_n net19 AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=1
XM99 net14 net15 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=2
XM101 net16 bias_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=2
XM102 net15 net15 net14 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=6
XM103 casc_p casc_p net14 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=4
XM104 casc_p casc_n net16 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM105 net15 casc_n net20 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM106 net17 bias_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=2
XM107 net6 casc_n net17 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM96 net18 bias_n net22 AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=1
XM108 net23 casc_n net18 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM109 bias_var_p casc_p net7 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM57 net19 bias_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=1
XM112 net20 casc_n net21 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM113 net22 bias_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=1
XM114 bias_var_p casc_n net23 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM115 Vx_hyst_n casc_n net12 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=3
XM118 net28 hyst0b_hv AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=6
XM119 net27 bias_p net28 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=6
XM120 Vx_hyst_p casc_p net27 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=6
XM121 net25 hyst1b_hv AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=16
XM122 net26 bias_p net25 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=18
XM123 Vx_hyst_p casc_p net26 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=18
XM124 Vfold_bot_p Voutb Vx_hyst_p AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=8
XM125 Vfold_bot_m Vout_int Vx_hyst_p AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=8
XM35 res_n_top res_n_top AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=4 nf=1 m=1
XM37 net31 bias_n net30 AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=4
XM41 net32 bias_n net33 AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=2
XM42 net30 trim1_hv AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=4
XM43 net33 trim0_hv AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=2
XM46 res_n_bot casc_n net31 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM47 res_n_bot casc_n net32 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM50 net35 trim2_hv res_n_top AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=16 nf=4 m=1
XM51 net34 trim2b_hv res_n_top AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=16 nf=4 m=1
XM52 net34 trim2_hv res_n_bot AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=16 nf=4 m=1
XM55 net35 trim2b_hv res_n_bot AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=16 nf=4 m=1
XM56 net36 bias_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=1
XM64 res_n_top casc_n net36 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM65 net37 trim0_hv res_n_top AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=16 nf=4 m=1
XM66 res_n_bot trim1_hv net37 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=16 nf=4 m=1
XR1 res_n_bot res_n_top AGND sky130_fd_pr__res_high_po_2p85 L=2.85*56 mult=1 m=1
XM71 net41 trim3b_hv AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=2
XM72 net40 bias_p net41 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=4
XM74 res_p_top casc_p net40 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM80 net38 trim4b_hv AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=4
XM81 net39 bias_p net38 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=8
XM82 res_p_top casc_p net39 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=8
XM83 Vfold_bot_m net46 net44 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1.5 W=8 nf=1 m=4
XM126 Vfold_bot_p net45 net44 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1.5 W=8 nf=1 m=4
XM127 net42 bias_var_tailp AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=12
XM128 net44 casc_p net42 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=12
XM129 net43 bias_p AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=2
XM130 res_p_bot casc_p net43 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XR2 res_p_bot res_p_top AGND sky130_fd_pr__res_high_po_2p85 L=2.85*56 mult=1 m=1
XM131 res_p_bot res_p_bot AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=1
XM132 net45 trim5_hv res_p_top AGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=16 nf=4 m=1
XM87 net49 bias_var_p AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=4
XM98 bias_var_tailn bias_var_tailn AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=2
XM100 net46 trim5b_hv res_p_top AGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=16 nf=4 m=1
XM135 res_p_bot trim5b_hv net45 AGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=16 nf=4 m=1
XM133 res_p_bot trim5_hv net46 AGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=16 nf=4 m=1
XM137 net47 trim4b_hv res_p_bot AGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=16 nf=4 m=1
XM136 res_p_top trim3b_hv net47 AGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=16 nf=4 m=1
x3 AVDD trim4b_hv trim4_hv trim[4] AGND DVDD DGND level_shifter_up
x9 AVDD trim5b_hv trim5_hv trim[5] AGND DVDD DGND level_shifter_up
XM134 net56 casc_p net48 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM138 net57 casc_p net49 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM139 net51 bias_p AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=2
XM140 bias_var_tailp casc_p net50 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=4
XM141 net7 bias_p net51 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=2
Vmeas_var_tailp net56 bias_var_n 0
.save i(vmeas_var_tailp)
Vmeas_var_tailn net57 bias_var_tailn 0
.save i(vmeas_var_tailn)
XM77 net53 ibias net52 AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=1
XM78 net54 ibias net53 AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=1
XM79 ibias ibias net54 AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=1
XM58 Vout Voutb DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM59 Vout Voutb DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM110 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=1.5 W=8 nf=1 m=34
XM111 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1.5 W=8 nf=1 m=36
XM116 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=15
XM117 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=14
XM142 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=32
XM143 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=32
XR3 AGND AGND AGND sky130_fd_pr__res_high_po_2p85 L=2.85*11.2 mult=1 m=1
XM144 casc_n casc_n casc_n AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=11
XM145 net55 bias_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5 L=4 W=2 nf=1 m=1
XM146 bias_stg2 casc_n net55 AGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM147 bias_stg2 bias_stg2 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=2
XM148 casc_p casc_p casc_p AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=20
XM149 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=2 nf=1 m=12
XR5 AGND AGND AGND sky130_fd_pr__res_high_po_2p85 L=2.85*11.2 mult=1 m=1
XR7 AGND AGND AGND sky130_fd_pr__res_high_po_2p85 L=2.85*11.2 mult=1 m=1
XR8 AGND AGND AGND sky130_fd_pr__res_high_po_2p85 L=2.85*11.2 mult=1 m=1
* noconn trim0b_hv
* noconn trim1b_hv
* noconn trim3_hv
* noconn trim4_hv
.ends


* expanding   symbol:  sky130_am_ip__ldo_01v8.sym # of pins=8
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_am_ip__ldo_01v8/xschem/sky130_am_ip__ldo_01v8.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_am_ip__ldo_01v8/xschem/sky130_am_ip__ldo_01v8.sch
.subckt sky130_am_ip__ldo_01v8 AVDD VOUT AVSS ENA VREF_EXT SEL_EXT DVDD DVSS
*.PININFO ENA:I AVDD:I AVSS:I VOUT:O SEL_EXT:I VREF_EXT:I DVDD:I DVSS:I
XM46 VX VBIAS_P AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=7 W=1 nf=1 m=1
XM48 net2 net2 AVSS AVSS sky130_fd_pr__nfet_g5v0d10v5 L=7 W=1 nf=1 m=1
XM52 VX VREF net1 AVSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM53 VY VM net1 AVSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM54 net1 VBIAS_N AVSS AVSS sky130_fd_pr__nfet_g5v0d10v5 L=9 W=3 nf=1 m=1
XM55 VERR net2 AVSS AVSS sky130_fd_pr__nfet_g5v0d10v5 L=7 W=1 nf=1 m=1
XM56 VY VBIAS_P AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=7 W=1 nf=1 m=1
XM57 VERR VBIAS_C VY AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM58 net2 VBIAS_C VX AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM59 AVSS VERR VPASS AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM60 VPASS VBIAS_P AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=7 W=1 nf=1 m=1
XR4 VM VOUT AVSS sky130_fd_pr__res_xhigh_po_0p35 L=180 mult=1 m=1
XR5 AVSS VM AVSS sky130_fd_pr__res_xhigh_po_0p35 L=360 mult=1 m=1
XM61 AVDD VPASS VOUT AVSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1000
XC1 VERR AVSS sky130_fd_pr__cap_mim_m3_1 W=15 L=15 m=3
XM62 net3 VBIAS_P AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=7 W=1 nf=1 m=1
XM63 VBIAS_P VBIAS_C net3 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM64 net4 VBIAS_P AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=7 W=1 nf=1 m=1
XM65 VBIAS_N VBIAS_C net4 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM66 VBIAS_P VBIAS_N net5 AVSS sky130_fd_pr__nfet_g5v0d10v5 L=9 W=1 nf=1 m=20
XM67 VBIAS_N VBIAS_N AVSS AVSS sky130_fd_pr__nfet_g5v0d10v5 L=9 W=1 nf=1 m=5
XM68 VBIAS_C VBIAS_C AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=10 W=1 nf=1 m=1
XM69 VBIAS_C VBIAS_N AVSS AVSS sky130_fd_pr__nfet_g5v0d10v5 L=9 W=1 nf=1 m=5
XM70 VDD_START VSTART VBIAS_N AVSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM71 net7 net7 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=1 nf=1 m=1
XM72 net6 net6 net7 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=1 nf=1 m=1
XM73 VSTART VSTART net6 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=1 nf=1 m=1
XM74 VSTART VBIAS_N AVSS AVSS sky130_fd_pr__nfet_g5v0d10v5 L=9 W=1 nf=1 m=5
XM75 NSEL_EXT sel_ext_3v3 AVSS AVSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM76 NSEL_EXT sel_ext_3v3 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2.5 nf=1 m=1
XM77 VREF NSEL_EXT VREF_INT AVSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM78 VREF sel_ext_3v3 VREF_EXT AVSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XC3 VREF AVSS sky130_fd_pr__cap_mim_m3_1 W=5 L=5 m=1
XR6 AVSS net5 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=40 mult=1 m=1
XM79 VREF_INT VBIAS_P AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=7 W=1 nf=1 m=1
XM80 net8 VREF_INT net9 AVSS sky130_fd_pr__nfet_g5v0d10v5 L=10 W=1 nf=1 m=1
XM81 VREF_INT VREF_INT net8 AVSS sky130_fd_pr__nfet_g5v0d10v5 L=10 W=1 nf=1 m=1
XM82 net9 VREF_INT AVSS AVSS sky130_fd_pr__nfet_g5v0d10v5 L=10 W=1 nf=1 m=1
XM83 NENA ena_3v3 AVSS AVSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM84 NENA ena_3v3 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2.5 nf=1 m=1
XM85 VBIAS_N NENA AVSS AVSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM86 VBIAS_C ena_3v3 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM87 VERR NENA AVSS AVSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM88 VBIAS_P ena_3v3 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM89 VPASS NENA AVSS AVSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM90 VDD_START NENA AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
x1 ENA DVDD DVSS DVSS AVDD AVDD ena_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x2 SEL_EXT DVDD DVSS DVSS AVDD AVDD sel_ext_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
.ends


* expanding   symbol:  sky130_ef_ip__cdac3v_12bit.sym # of pins=25
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/sky130_ef_ip__cdac3v_12bit.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/sky130_ef_ip__cdac3v_12bit.sch
.subckt sky130_ef_ip__cdac3v_12bit SELD0 SELD1 SELD2 SELD3 SELD4 SELD5 SELD6 SELD7 SELD8 SELD9 VDD DVDD DVSS VSS VH VL OUT RST
+ OUTNC SELD10 SELD11 VCM Vref VIN HOLD
*.PININFO SELD0:I SELD1:I SELD2:I SELD3:I SELD4:I SELD5:I SELD6:I SELD7:I SELD8:I SELD9:I VDD:B DVDD:B DVSS:B VH:B VL:B VSS:B
*+ RST:I OUT:O OUTNC:O SELD10:I SELD11:I VIN:B Vref:B VCM:B HOLD:I
x4 D8 D0 D4 OUTNC D9 D5 D1 OUT D2 D6 VSS D7 D3 D10 D11 Vref EF_BANK_CAP_12
x3 D0 sel0_3v3 D1 sel1_3v3 sel2_3v3 D2 sel3_3v3 sel4_3v3 D3 sel5_3v3 D4 sel6_3v3 sel7_3v3 D5 sel8_3v3 D6 sel9_3v3 D7 D8 D9 VDD
+ DVSS VH VL VSS D10 D11 sel10_3v3 sel11_3v3 VCM rst_3v3 EF_AMUX0201_ARRAY1
x1 OUTNC OUT VDD VSS hold_3v3 VIN DVSS holdb_3v3 EF_SW_RST
x2 SELD3 sel3_3v3 sel7_3v3 SELD7 sel11_3v3 SELD11 SELD6 sel6_3v3 SELD10 sel2_3v3 sel10_3v3 SELD2 sel1_3v3 sel5_3v3 SELD5 SELD1
+ SELD9 sel9_3v3 VDD DVSS sel0_3v3 SELD4 sel4_3v3 sel8_3v3 SELD8 DVDD SELD0 hold_3v3 HOLD rst_3v3 RST holdb_3v3 cdac_lvlshift_array
.ends


* expanding   symbol:  sky130_ef_ip__rheostat_8bit.sym # of pins=15
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rheostat_8bit/xschem/sky130_ef_ip__rheostat_8bit.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rheostat_8bit/xschem/sky130_ef_ip__rheostat_8bit.sch
.subckt sky130_ef_ip__rheostat_8bit dvdd vss dvss vdd b0 Vhigh b1 b2 b3 out b4 b5 b6 b7 Vlow
*.PININFO out:B vss:B vdd:B Vhigh:B Vlow:B b0:I b1:I b2:I b3:I b4:I b5:I b6:I b7:I dvdd:B dvss:B
x1 vdd vss b3a b4a b3b b4b b5a Vhigh b6a b0a net3 b6b b5b b0b b1a b1b b2a b2b net1 net6 net5 rheo_half
x2 vdd vss b3a b4a b3b b4b b5a net6 b6a b0a net5 b6b b5b b0b b1a b1b b2a b2b net2 Vlow net4 rheo_half
x3 vdd b7b out net1 b7a vss passtrans
x7 vdd dvdd b7a b7b b7 dvss rheo_level_shifter
x8 vdd dvdd b6a b6b b6 dvss rheo_level_shifter
x9 vdd dvdd b5a b5b b5 dvss rheo_level_shifter
x10 vdd dvdd b4a b4b b4 dvss rheo_level_shifter
x11 vdd dvdd b3a b3b b3 dvss rheo_level_shifter
x12 vdd dvdd b2a b2b b2 dvss rheo_level_shifter
x13 vdd dvdd b1a b1b b1 dvss rheo_level_shifter
x14 vdd dvdd b0a b0b b0 dvss rheo_level_shifter
x15 vdd b7a out net2 b7b vss passtrans
x18 vdd net4 Vlow net7 vss net8 rheo_column_dummy
x5 vdd net8 net7 net9 vss net9 rheo_column_dummy
x4 vdd net10 net11 Vhigh vss net3 rheo_column_dummy
x16 vdd net12 net12 net11 vss net10 rheo_column_dummy
.ends


* expanding   symbol:  sky130_icrg_ip__ulpcomp2.sym # of pins=9
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_icrg_ip__ulpcomp/xschem/sky130_icrg_ip__ulpcomp2.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_icrg_ip__ulpcomp/xschem/sky130_icrg_ip__ulpcomp2.sch
.subckt sky130_icrg_ip__ulpcomp2 dvdd avdd ena vout vinn vinp clk dvss avss
*.PININFO avdd:I vinp:I vinn:I vout:O dvdd:I clk:I ena:I dvss:I avss:I
x1 dvddb clka clk clkb dvss Stage0_clk_inv
x2 avdd enab clka vinn vinp net2 net1 avss dvss dvdd Stage1
x3 dvdd enab dvddb clkb vout net2 net1 dvss Stage2_latch
x4 dvdd ena enab dvss Stage0_ena_inv
.ends


* expanding   symbol:  sky130_od_ip__tempsensor_ext_vp.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_od_ip__tempsensor/xschem/sky130_od_ip__tempsensor_ext_vp.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_od_ip__tempsensor/xschem/sky130_od_ip__tempsensor_ext_vp.sch
.subckt sky130_od_ip__tempsensor_ext_vp vbe1_out vdd vss vbg ena vbe2_out
*.PININFO vdd:I vss:I vbe2_out:O vbe1_out:O ena:I vbg:I
XQ_BL1 vss vss vbe1 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XQ_BR1 vss vss vbe2 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XM4 net2 vbg net1 vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM5 vp vp net1 vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM7 vp net2 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XM8 net2 net2 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XM3 vp ena vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XM6 net1 ena vss vss sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
x1 vdd vss ena vbe1 vbe1_out buffer
x2 vdd vss ena vbe2 vbe2_out buffer
XM1 vbe1 vp vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XM2 vbe2 vp vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=5
XD1 vss ena sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
XD2 vss vbg sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
.ends


* expanding   symbol:  sky130_vbl_ip__overvoltage.sym # of pins=12
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_vbl_ip__overvoltage/xschem/sky130_vbl_ip__overvoltage.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_vbl_ip__overvoltage/xschem/sky130_vbl_ip__overvoltage.sch
.subckt sky130_vbl_ip__overvoltage ovout vtrip[0] dvss avss avdd dvdd ibias vbg ena vtrip[3] vtrip[2] vtrip[1]
*.PININFO avdd:B dvdd:B ena:I avss:B vtrip[3]:I ovout:O vbg:I vtrip[2]:I vtrip[1]:I vtrip[0]:I ibias:I dvss:B
x1 dvdd ovout vbg net17 ena ibias dvss comp_hyst
x2 net2 net3 net4 net5 net6 net7 net8 avdd avss net9 A NotA B NotB C net17 NotC D NotD net1 net10 net11 net12 net13 net14 net15
+ net16 ov_multiplexer
x3 avdd net2 net3 net4 net5 net6 net7 net8 net9 net1 net10 net11 net12 net13 net14 net15 net16 avss ena ov_voltage_divider
x4 avdd dvdd vtrip[3] A NotA avss dvss ov_level_shifter
x5 avdd dvdd vtrip[2] B NotB avss dvss ov_level_shifter
x6 avdd dvdd vtrip[1] C NotC avss dvss ov_level_shifter
x7 avdd dvdd vtrip[0] D NotD avss dvss ov_level_shifter
.ends


* expanding   symbol:  sky130_ef_ip__rdac3v_8bit.sym # of pins=16
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rdac3v_8bit/xschem/sky130_ef_ip__rdac3v_8bit.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rdac3v_8bit/xschem/sky130_ef_ip__rdac3v_8bit.sch
.subckt sky130_ef_ip__rdac3v_8bit dvdd vss dvss vdd b0 Vhigh b1 b2 b3 out b4 b5 ena b6 b7 Vlow
*.PININFO out:O vss:B vdd:B Vhigh:B Vlow:B ena:I b0:I b1:I b2:I b3:I b4:I b5:I b6:I b7:I dvdd:B dvss:B
x1 vdd vss b3a b4a b3b b4b b5a Vhigh b6a b0a net3 b6b b5b b0b b1a b1b b2a b2b net1 net6 net5 dac_half
x2 vdd vss b3a b4a b3b b4b b5a net6 b6a b0a net5 b6b b5b b0b b1a b1b b2a b2b net2 Vlow net4 dac_half
x3 vdd b7b out_unbuf net1 b7a vss passtrans
x7 vdd dvdd b7a b7b b7 dvss level_shifter
x8 vdd dvdd b6a b6b b6 dvss level_shifter
x9 vdd dvdd b5a b5b b5 dvss level_shifter
x10 vdd dvdd b4a b4b b4 dvss level_shifter
x11 vdd dvdd b3a b3b b3 dvss level_shifter
x12 vdd dvdd b2a b2b b2 dvss level_shifter
x13 vdd dvdd b1a b1b b1 dvss level_shifter
x14 vdd dvdd b0a b0b b0 dvss level_shifter
x15 vdd b7a out_unbuf net2 b7b vss passtrans
x18 vdd net4 Vlow net7 vss net8 dac_column_dummy
x5 vdd net8 net7 net9 vss net9 dac_column_dummy
x4 vdd net10 net11 Vhigh vss net3 dac_column_dummy
x16 vdd net12 net12 net11 vss net10 dac_column_dummy
x6 vdd out ena vss out_unbuf dvss follower_amp
.ends


* expanding   symbol:  switch_array_18.sym # of pins=34
** sym_path: /home/tim/gits/frigate_analog/xschem/switch_array_18.sym
** sch_path: /home/tim/gits/frigate_analog/xschem/switch_array_18.sch
.subckt switch_array_18 avdd dvdd dvss avss adc1 comp_n ulpcomp_n right_instramp_to_ulpcomp_n[1] right_instramp_to_ulpcomp_n[0]
+ right_instramp_out right_hgbw_opamp_to_ulpcomp_n[1] right_hgbw_opamp_to_ulpcomp_n[0] right_lp_opamp_to_ulpcomp_p[1] right_lp_opamp_to_ulpcomp_p[0]
+ left_lp_opamp_to_ulpcomp_n[1] left_lp_opamp_to_ulpcomp_n[0] left_hgbw_opamp_to_ulpcomp_p[1] left_hgbw_opamp_to_ulpcomp_p[0] left_instramp_to_ulpcomp_p[1]
+ left_instramp_to_ulpcomp_p[0] right_hgbw_opamp_out right_instramp_to_comp_n[1] right_instramp_to_comp_n[0] right_hgbw_opamp_to_comp_n[1]
+ right_hgbw_opamp_to_comp_n[0] right_lp_opamp_to_comp_p[1] right_lp_opamp_to_comp_p[0] left_lp_opamp_to_comp_n[1] left_lp_opamp_to_comp_n[0]
+ left_hgbw_opamp_to_comp_p[1] left_hgbw_opamp_to_comp_p[0] left_instramp_to_comp_p[1] left_instramp_to_comp_p[0] right_lp_opamp_out right_instramp_to_adc1[1]
+ right_instramp_to_adc1[0] right_hgbw_opamp_to_adc1[1] right_hgbw_opamp_to_adc1[0] right_lp_opamp_to_adc0[1] right_lp_opamp_to_adc0[0]
+ left_lp_opamp_to_adc1[1] left_lp_opamp_to_adc1[0] left_hgbw_opamp_to_adc0[1] left_hgbw_opamp_to_adc0[0] left_lp_opamp_out left_instramp_to_adc0[1]
+ left_instramp_to_adc0[0] left_hgbw_opamp_out left_instramp_out adc0 ulpcomp_p comp_p
*.PININFO right_instramp_out:B right_hgbw_opamp_out:B left_lp_opamp_out:B right_lp_opamp_out:B left_hgbw_opamp_out:B
*+ left_instramp_out:B ulpcomp_n:B comp_n:B adc1:B comp_p:B ulpcomp_p:B adc0:B avdd:B dvdd:B dvss:B avss:B right_instramp_to_ulpcomp_n[1:0]:I
*+ right_hgbw_opamp_to_ulpcomp_n[1:0]:I right_lp_opamp_to_ulpcomp_p[1:0]:I left_lp_opamp_to_ulpcomp_n[1:0]:I right_instramp_to_comp_n[1:0]:I
*+ right_instramp_to_adc1[1:0]:I left_hgbw_opamp_to_ulpcomp_p[1:0]:I left_instramp_to_ulpcomp_p[1:0]:I right_hgbw_opamp_to_comp_n[1:0]:I
*+ right_lp_opamp_to_comp_p[1:0]:I left_lp_opamp_to_comp_n[1:0]:I left_hgbw_opamp_to_comp_p[1:0]:I left_instramp_to_comp_p[1:0]:I right_hgbw_opamp_to_adc1[1:0]:I
*+ right_lp_opamp_to_adc0[1:0]:I left_lp_opamp_to_adc1[1:0]:I left_hgbw_opamp_to_adc0[1:0]:I left_instramp_to_adc0[1:0]:I
x4 avss right_instramp_to_ulpcomp_n[0] right_instramp_out ulpcomp_n avdd dvdd dvss right_instramp_to_ulpcomp_n[1]
+ isolated_switch_large
x5 avss right_hgbw_opamp_to_ulpcomp_n[0] right_hgbw_opamp_out ulpcomp_n avdd dvdd dvss right_hgbw_opamp_to_ulpcomp_n[1]
+ isolated_switch_large
x6 avss left_lp_opamp_to_ulpcomp_n[0] left_lp_opamp_out ulpcomp_n avdd dvdd dvss left_lp_opamp_to_ulpcomp_n[1]
+ isolated_switch_large
x7 avss right_lp_opamp_to_comp_p[0] right_lp_opamp_out comp_p avdd dvdd dvss right_lp_opamp_to_comp_p[1] isolated_switch_large
x8 avss left_hgbw_opamp_to_comp_p[0] left_hgbw_opamp_out comp_p avdd dvdd dvss left_hgbw_opamp_to_comp_p[1] isolated_switch_large
x9 avss left_instramp_to_comp_p[0] left_instramp_out comp_p avdd dvdd dvss left_instramp_to_comp_p[1] isolated_switch_large
x10 avss right_lp_opamp_to_adc0[0] right_lp_opamp_out adc0 avdd dvdd dvss right_lp_opamp_to_adc0[1] isolated_switch_large
x11 avss left_hgbw_opamp_to_adc0[0] left_hgbw_opamp_out adc0 avdd dvdd dvss left_hgbw_opamp_to_adc0[1] isolated_switch_large
x12 avss left_instramp_to_adc0[0] left_instramp_out adc0 avdd dvdd dvss left_instramp_to_adc0[1] isolated_switch_large
x1 avss right_instramp_to_comp_n[0] right_instramp_out comp_n avdd dvdd dvss right_instramp_to_comp_n[1] isolated_switch_large
x2 avss right_hgbw_opamp_to_comp_n[0] right_hgbw_opamp_out comp_n avdd dvdd dvss right_hgbw_opamp_to_comp_n[1]
+ isolated_switch_large
x3 avss left_lp_opamp_to_comp_n[0] left_lp_opamp_out comp_n avdd dvdd dvss left_lp_opamp_to_comp_n[1] isolated_switch_large
x13 avss right_lp_opamp_to_ulpcomp_p[0] right_lp_opamp_out ulpcomp_p avdd dvdd dvss right_lp_opamp_to_ulpcomp_p[1]
+ isolated_switch_large
x14 avss left_hgbw_opamp_to_ulpcomp_p[0] left_hgbw_opamp_out ulpcomp_p avdd dvdd dvss left_hgbw_opamp_to_ulpcomp_p[1]
+ isolated_switch_large
x15 avss left_instramp_to_ulpcomp_p[0] left_instramp_out ulpcomp_p avdd dvdd dvss left_instramp_to_ulpcomp_p[1]
+ isolated_switch_large
x16 avss right_instramp_to_adc1[0] right_instramp_out adc1 avdd dvdd dvss right_instramp_to_adc1[1] isolated_switch_large
x17 avss right_hgbw_opamp_to_adc1[0] right_hgbw_opamp_out adc1 avdd dvdd dvss right_hgbw_opamp_to_adc1[1] isolated_switch_large
x18 avss left_lp_opamp_to_adc1[0] left_lp_opamp_out adc1 avdd dvdd dvss left_lp_opamp_to_adc1[1] isolated_switch_large
.ends


* expanding   symbol:  switch_array_14.sym # of pins=30
** sym_path: /home/tim/gits/frigate_analog/xschem/switch_array_14.sym
** sch_path: /home/tim/gits/frigate_analog/xschem/switch_array_14.sch
.subckt switch_array_14 avdd dvdd dvss avss right_instramp_to_amuxbusA[1] right_instramp_to_amuxbusA[0] right_instramp_out
+ left_hgbw_opamp_to_amuxbusB[1] left_hgbw_opamp_to_amuxbusB[0] left_lp_opamp_to_amuxbusA[1] left_lp_opamp_to_amuxbusA[0] right_lp_opamp_to_amuxbusB[1]
+ right_lp_opamp_to_amuxbusB[0] right_hgbw_opamp_to_amuxbusA[1] right_hgbw_opamp_to_amuxbusA[0] left_instramp_to_amuxbusB[1] left_instramp_to_amuxbusB[0]
+ right_hgbw_opamp_out right_instramp_to_analog0[1] right_instramp_to_analog0[0] left_hgbw_opamp_to_analog1[1] left_hgbw_opamp_to_analog1[0]
+ left_lp_opamp_to_analog0[1] left_lp_opamp_to_analog0[0] right_lp_opamp_to_analog1[1] right_lp_opamp_to_analog1[0] right_hgbw_opamp_to_analog0[1]
+ right_hgbw_opamp_to_analog0[0] left_instramp_to_analog1[1] left_instramp_to_analog1[0] right_lp_opamp_out left_lp_opamp_out left_hgbw_opamp_out
+ left_instramp_out analog1 analog1_core analog0 analog0_core amuxbusB amuxbusA analog1_connect[1] analog1_connect[0] analog0_connect[1]
+ analog0_connect[0]
*.PININFO right_instramp_out:B right_hgbw_opamp_out:B right_lp_opamp_out:B left_lp_opamp_out:B left_hgbw_opamp_out:B
*+ left_instramp_out:B analog0_core:B avdd:B dvdd:B dvss:B avss:B right_instramp_to_analog0[1:0]:I left_hgbw_opamp_to_analog1[1:0]:I
*+ left_lp_opamp_to_analog0[1:0]:I right_lp_opamp_to_analog1[1:0]:I right_instramp_to_amuxbusA[1:0]:I right_hgbw_opamp_to_analog0[1:0]:I
*+ left_instramp_to_analog1[1:0]:I left_hgbw_opamp_to_amuxbusB[1:0]:I left_lp_opamp_to_amuxbusA[1:0]:I right_lp_opamp_to_amuxbusB[1:0]:I
*+ right_hgbw_opamp_to_amuxbusA[1:0]:I left_instramp_to_amuxbusB[1:0]:I analog0:B analog1_core:B analog1:B amuxbusA:B amuxbusB:B analog1_connect[1:0]:I
*+ analog0_connect[1:0]:I
x10 avss analog1_connect[0] analog1 analog1_core avdd dvdd dvss analog1_connect[1] isolated_switch_xlarge
x11 avss analog0_connect[0] analog0 analog0_core avdd dvdd dvss analog0_connect[1] isolated_switch_xlarge
x1 avss left_instramp_to_amuxbusB[0] left_instramp_out amuxbusB avdd dvdd dvss left_instramp_to_amuxbusB[1] isolated_switch_xlarge
x2 avss left_hgbw_opamp_to_amuxbusB[0] left_hgbw_opamp_out amuxbusB avdd dvdd dvss left_hgbw_opamp_to_amuxbusB[1]
+ isolated_switch_xlarge
x3 avss right_lp_opamp_to_amuxbusB[0] right_lp_opamp_out amuxbusB avdd dvdd dvss right_lp_opamp_to_amuxbusB[1]
+ isolated_switch_xlarge
x4 avss right_lp_opamp_to_analog1[0] right_lp_opamp_out analog1_core avdd dvdd dvss right_lp_opamp_to_analog1[1]
+ isolated_switch_xlarge
x5 avss left_hgbw_opamp_to_analog1[0] left_hgbw_opamp_out analog1_core avdd dvdd dvss left_hgbw_opamp_to_analog1[1]
+ isolated_switch_xlarge
x6 avss left_instramp_to_analog1[0] left_instramp_out analog1_core avdd dvdd dvss left_instramp_to_analog1[1]
+ isolated_switch_xlarge
x7 avss right_instramp_to_analog0[0] right_instramp_out analog0_core avdd dvdd dvss right_instramp_to_analog0[1]
+ isolated_switch_xlarge
x8 avss right_hgbw_opamp_to_analog0[0] right_hgbw_opamp_out analog0_core avdd dvdd dvss right_hgbw_opamp_to_analog0[1]
+ isolated_switch_xlarge
x9 avss left_lp_opamp_to_analog0[0] left_lp_opamp_out analog0_core avdd dvdd dvss left_lp_opamp_to_analog0[1]
+ isolated_switch_xlarge
x12 avss left_lp_opamp_to_amuxbusA[0] left_lp_opamp_out amuxbusA avdd dvdd dvss left_lp_opamp_to_amuxbusA[1]
+ isolated_switch_xlarge
x13 avss right_hgbw_opamp_to_amuxbusA[0] right_hgbw_opamp_out amuxbusA avdd dvdd dvss right_hgbw_opamp_to_amuxbusA[1]
+ isolated_switch_xlarge
x14 avss right_instramp_to_amuxbusA[0] right_instramp_out amuxbusA avdd dvdd dvss right_instramp_to_amuxbusA[1]
+ isolated_switch_xlarge
.ends


* expanding   symbol:  switch_array_4.sym # of pins=16
** sym_path: /home/tim/gits/frigate_analog/xschem/switch_array_4.sym
** sch_path: /home/tim/gits/frigate_analog/xschem/switch_array_4.sch
.subckt switch_array_4 avdd dvdd dvss avss channel0_out channel0_in_to_out[1] channel0_in_to_out[0] channel0_in
+ channel1_in_to_out[1] channel1_in_to_out[0] channel2_in_to_out[1] channel2_in_to_out[0] channel3_in_to_out[1] channel3_in_to_out[0] channel1_out
+ channel1_in channel2_out channel2_in channel3_out channel3_in
*.PININFO channel0_in:B avdd:B dvdd:B dvss:B avss:B channel0_in_to_out[1:0]:I channel0_out:B channel1_in:B channel1_out:B
*+ channel2_in:B channel2_out:B channel3_in:B channel3_out:B channel1_in_to_out[1:0]:I channel2_in_to_out[1:0]:I channel3_in_to_out[1:0]:I
x1 avss channel0_in_to_out[0] channel0_out channel0_in avdd dvdd dvss channel0_in_to_out[1] isolated_switch_xlarge
x2 avss channel1_in_to_out[0] channel1_out channel1_in avdd dvdd dvss channel1_in_to_out[1] isolated_switch_xlarge
x3 avss channel2_in_to_out[0] channel2_out channel2_in avdd dvdd dvss channel2_in_to_out[1] isolated_switch_xlarge
x4 avss channel3_in_to_out[0] channel3_out channel3_in avdd dvdd dvss channel3_in_to_out[1] isolated_switch_xlarge
.ends


* expanding   symbol:  simple_switch_array_32.sym # of pins=60
** sym_path: /home/tim/gits/frigate_analog/xschem/simple_switch_array_32.sym
** sch_path: /home/tim/gits/frigate_analog/xschem/simple_switch_array_32.sch
.subckt simple_switch_array_32 vdda0 vssa0 vccd0 vssd0 analog1 amuxbusA amuxbusB analog0 right_instramp_n_to_analog1
+ right_instramp_p_to_amuxbusA right_instramp_n_to_amuxbusB right_instramp_p_to_analog0 right_instramp_n right_hgbw_opamp_n_to_analog1 right_instramp_p
+ right_hgbw_opamp_n_to_amuxbusB right_hgbw_opamp_p_to_amuxbusA right_hgbw_opamp_p_to_analog0 right_hgbw_opamp_n right_hgbw_opamp_p right_lp_opamp_n
+ right_lp_opamp_p right_lp_opamp_n_to_analog1 right_lp_opamp_p_to_amuxbusA right_lp_opamp_p_to_analog0 right_lp_opamp_n_to_amuxbusB left_instramp_n
+ left_instramp_p left_hgbw_opamp_n left_hgbw_opamp_p left_lp_opamp_n_to_analog1 left_lp_opamp_p_to_amuxbusA left_lp_opamp_n_to_amuxbusB
+ left_lp_opamp_p_to_analog0 left_lp_opamp_n left_lp_opamp_p ulpcomp_p ulpcomp_n left_hgbw_opamp_n_to_analog1 left_hgbw_opamp_p_to_analog0
+ left_hgbw_opamp_n_to_amuxbusB left_hgbw_opamp_p_to_amuxbusA comp_p comp_n adc0 adc1 left_instramp_n_to_analog1 dac0 left_instramp_p_to_analog0
+ left_instramp_n_to_amuxbusB left_instramp_p_to_amuxbusA dac1 ulpcomp_p_to_analog1 ulpcomp_n_to_analog0 comp_p_to_analog1 comp_n_to_analog0 adc0_to_analog1
+ adc1_to_analog0 dac0_to_analog1 dac1_to_analog0
*.PININFO vccd0:B right_instramp_n_to_analog1:I vdda0:B vssa0:B vssd0:B right_hgbw_opamp_n_to_analog1:I
*+ right_lp_opamp_n_to_analog1:I left_lp_opamp_n_to_analog1:I left_hgbw_opamp_n_to_analog1:I left_instramp_n_to_analog1:I ulpcomp_p_to_analog1:I
*+ comp_p_to_analog1:I adc0_to_analog1:I dac0_to_analog1:I analog1:B right_instramp_p_to_analog0:I right_hgbw_opamp_p_to_analog0:I
*+ right_lp_opamp_p_to_analog0:I left_lp_opamp_p_to_analog0:I left_hgbw_opamp_p_to_analog0:I left_instramp_p_to_analog0:I ulpcomp_n_to_analog0:I
*+ comp_n_to_analog0:I adc1_to_analog0:I dac1_to_analog0:I analog0:B amuxbusA:B right_instramp_p_to_amuxbusA:I right_hgbw_opamp_p_to_amuxbusA:I
*+ right_lp_opamp_p_to_amuxbusA:I left_lp_opamp_p_to_amuxbusA:I left_hgbw_opamp_p_to_amuxbusA:I left_instramp_p_to_amuxbusA:I amuxbusB:B
*+ right_instramp_n_to_amuxbusB:I right_hgbw_opamp_n_to_amuxbusB:I right_lp_opamp_n_to_amuxbusB:I left_lp_opamp_n_to_amuxbusB:I left_hgbw_opamp_n_to_amuxbusB:I
*+ left_instramp_n_to_amuxbusB:I right_instramp_n:B right_instramp_p:B right_hgbw_opamp_n:B right_hgbw_opamp_p:B right_lp_opamp_n:B right_lp_opamp_p:B
*+ left_instramp_n:B left_instramp_p:B left_hgbw_opamp_n:B left_hgbw_opamp_p:B left_lp_opamp_n:B left_lp_opamp_p:B ulpcomp_p:B ulpcomp_n:B comp_p:B
*+ comp_n:B adc0:B adc1:B dac0:B dac1:B
x1 vssa0 right_instramp_n_to_analog1 analog1 right_instramp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x2 vssa0 right_hgbw_opamp_n_to_analog1 analog1 right_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x3 vssa0 right_lp_opamp_n_to_analog1 analog1 right_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x4 vssa0 left_lp_opamp_n_to_analog1 analog1 left_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x5 vssa0 left_hgbw_opamp_n_to_analog1 analog1 left_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x6 vssa0 left_instramp_n_to_analog1 analog1 left_instramp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x7 vssa0 ulpcomp_p_to_analog1 analog1 ulpcomp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x8 vssa0 comp_p_to_analog1 analog1 comp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x9 vssa0 adc0_to_analog1 analog1 adc0 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x10 vssa0 dac0_to_analog1 analog1 dac0 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x11 vssa0 right_instramp_p_to_analog0 analog0 right_instramp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x12 vssa0 right_hgbw_opamp_p_to_analog0 analog0 right_hgbw_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x13 vssa0 right_lp_opamp_p_to_analog0 analog0 right_lp_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x14 vssa0 left_lp_opamp_p_to_analog0 analog0 left_lp_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x15 vssa0 left_hgbw_opamp_p_to_analog0 analog0 left_hgbw_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x16 vssa0 left_instramp_p_to_analog0 analog0 left_instramp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x17 vssa0 ulpcomp_n_to_analog0 analog0 ulpcomp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x18 vssa0 comp_n_to_analog0 analog0 comp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x19 vssa0 adc1_to_analog0 analog0 adc1 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x20 vssa0 dac1_to_analog0 analog0 dac1 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x21 vssa0 right_instramp_n_to_amuxbusB amuxbusB right_instramp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x22 vssa0 right_hgbw_opamp_n_to_amuxbusB amuxbusB right_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x23 vssa0 right_lp_opamp_n_to_amuxbusB amuxbusB right_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x24 vssa0 left_lp_opamp_n_to_amuxbusB amuxbusB left_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x25 vssa0 left_hgbw_opamp_n_to_amuxbusB amuxbusB left_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x26 vssa0 left_instramp_n_to_amuxbusB amuxbusB left_instramp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x28 vssa0 right_instramp_p_to_amuxbusA amuxbusA right_instramp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x29 vssa0 right_hgbw_opamp_p_to_amuxbusA amuxbusA right_hgbw_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x30 vssa0 right_lp_opamp_p_to_amuxbusA amuxbusA right_lp_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x31 vssa0 left_lp_opamp_p_to_amuxbusA amuxbusA left_lp_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x32 vssa0 left_hgbw_opamp_p_to_amuxbusA amuxbusA left_hgbw_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x33 vssa0 left_instramp_p_to_amuxbusA amuxbusA left_instramp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
.ends


* expanding   symbol:  simple_switch_array_53.sym # of pins=82
** sym_path: /home/tim/gits/frigate_analog/xschem/simple_switch_array_53.sym
** sch_path: /home/tim/gits/frigate_analog/xschem/simple_switch_array_53.sch
.subckt simple_switch_array_53 vdda0 vssa0 vccd0 vssd0 vbgtc vbgsc left_vref tempsense right_vref voutref vinref
+ right_instramp_p_to_left_vref right_instramp_n_to_right_vref right_instramp_p_to_tempsense right_instramp_n_to_vinref right_instramp_p_to_voutref
+ right_instramp_n right_instramp_p right_hgbw_opamp_n_to_vbgsc right_hgbw_opamp_n right_hgbw_opamp_p right_hgbw_opamp_n_to_right_vref
+ right_hgbw_opamp_p_to_left_vref right_hgbw_opamp_n_to_vinref right_hgbw_opamp_p_to_voutref right_lp_opamp_n right_lp_opamp_p right_lp_opamp_n_to_vbgtc
+ left_instramp_n left_instramp_p right_lp_opamp_n_to_right_vref right_lp_opamp_p_to_left_vref right_lp_opamp_p_to_voutref
+ right_lp_opamp_n_to_vinref left_hgbw_opamp_n left_lp_opamp_n_to_vbgsc left_hgbw_opamp_p left_lp_opamp_n left_lp_opamp_p right_lp_opamp_p_to_tempsense
+ left_lp_opamp_n_to_right_vref left_lp_opamp_p_to_left_vref left_lp_opamp_p_to_voutref left_lp_opamp_n_to_vinref ulpcomp_p ulpcomp_n
+ left_hgbw_opamp_p_to_tempsense comp_p comp_n left_hgbw_opamp_n_to_right_vref left_hgbw_opamp_p_to_left_vref left_hgbw_opamp_p_to_voutref
+ left_hgbw_opamp_n_to_vinref adc0 adc1 left_instramp_n_to_right_vref left_instramp_p_to_tempsense left_instramp_p_to_left_vref left_instramp_p_to_voutref
+ left_instramp_n_to_vinref ulpcomp_p_to_vbgtc ulpcomp_n_to_vbgsc ulpcomp_n_to_vinref ulpcomp_p_to_left_vref ulpcomp_n_to_right_vref ulpcomp_p_to_tempsense
+ ulpcomp_p_to_voutref comp_p_to_vbgtc comp_n_to_vbgsc comp_n_to_vinref comp_p_to_left_vref comp_n_to_right_vref comp_p_to_tempsense comp_p_to_voutref
+ adc0_to_vbgtc adc1_to_vbgsc adc1_to_vinref adc1_to_right_vref adc0_to_left_vref adc0_to_tempsense adc0_to_voutref left_hgbw_opamp_n_to_vbgtc
*.PININFO vccd0:B vdda0:B vssa0:B vssd0:B left_hgbw_opamp_n_to_vbgtc:I right_lp_opamp_n_to_vbgtc:I ulpcomp_p_to_vbgtc:I
*+ comp_p_to_vbgtc:I adc0_to_vbgtc:I vbgtc:B left_lp_opamp_n_to_vbgsc:I right_hgbw_opamp_n_to_vbgsc:I ulpcomp_n_to_vbgsc:I comp_n_to_vbgsc:I
*+ adc1_to_vbgsc:I vbgsc:B right_vref:B left_instramp_p_to_tempsense:I left_hgbw_opamp_p_to_tempsense:I right_lp_opamp_p_to_tempsense:I
*+ right_instramp_p_to_tempsense:I tempsense:B right_instramp_n_to_right_vref:I right_hgbw_opamp_n_to_right_vref:I right_lp_opamp_n_to_right_vref:I
*+ left_lp_opamp_n_to_right_vref:I left_hgbw_opamp_n_to_right_vref:I left_instramp_n_to_right_vref:I right_instramp_n:B right_instramp_p:B right_hgbw_opamp_n:B
*+ right_hgbw_opamp_p:B right_lp_opamp_n:B right_lp_opamp_p:B left_instramp_n:B left_instramp_p:B left_hgbw_opamp_n:B left_hgbw_opamp_p:B
*+ left_lp_opamp_n:B left_lp_opamp_p:B ulpcomp_p:B ulpcomp_n:B comp_p:B comp_n:B adc0:B adc1:B ulpcomp_p_to_tempsense:I comp_p_to_tempsense:I
*+ adc0_to_tempsense:I ulpcomp_n_to_right_vref:I comp_n_to_right_vref:I adc1_to_right_vref:I ulpcomp_p_to_left_vref:I comp_p_to_left_vref:I
*+ adc0_to_left_vref:I ulpcomp_n_to_vinref:I comp_n_to_vinref:I adc1_to_vinref:I ulpcomp_p_to_voutref:I comp_p_to_voutref:I adc0_to_voutref:I
*+ left_vref:B right_instramp_p_to_left_vref:I right_hgbw_opamp_p_to_left_vref:I right_lp_opamp_p_to_left_vref:I left_lp_opamp_p_to_left_vref:I
*+ left_hgbw_opamp_p_to_left_vref:I left_instramp_p_to_left_vref:I vinref:B right_instramp_n_to_vinref:I right_hgbw_opamp_n_to_vinref:I right_lp_opamp_n_to_vinref:I
*+ left_lp_opamp_n_to_vinref:I left_hgbw_opamp_n_to_vinref:I left_instramp_n_to_vinref:I voutref:B right_instramp_p_to_voutref:I right_hgbw_opamp_p_to_voutref:I
*+ right_lp_opamp_p_to_voutref:I left_lp_opamp_p_to_voutref:I left_hgbw_opamp_p_to_voutref:I left_instramp_p_to_voutref:I
x2 vssa0 left_hgbw_opamp_n_to_vbgtc vbgtc left_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x4 vssa0 right_lp_opamp_n_to_vbgtc vbgtc right_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x7 vssa0 ulpcomp_p_to_vbgtc vbgtc ulpcomp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x8 vssa0 comp_p_to_vbgtc vbgtc comp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x9 vssa0 adc0_to_vbgtc vbgtc adc0 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x13 vssa0 left_lp_opamp_n_to_vbgsc vbgsc left_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x15 vssa0 right_hgbw_opamp_n_to_vbgsc vbgsc right_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x17 vssa0 ulpcomp_n_to_vbgsc vbgsc ulpcomp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x18 vssa0 comp_n_to_vbgsc vbgsc comp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x19 vssa0 adc1_to_vbgsc vbgsc adc1 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x21 vssa0 right_instramp_n_to_right_vref right_vref right_instramp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x22 vssa0 right_hgbw_opamp_n_to_right_vref right_vref right_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x23 vssa0 right_lp_opamp_n_to_right_vref right_vref right_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x24 vssa0 left_lp_opamp_n_to_right_vref right_vref left_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x25 vssa0 left_hgbw_opamp_n_to_right_vref right_vref left_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x26 vssa0 left_instramp_n_to_right_vref right_vref left_instramp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x28 vssa0 left_instramp_p_to_tempsense tempsense left_instramp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x29 vssa0 left_hgbw_opamp_p_to_tempsense tempsense left_hgbw_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x31 vssa0 right_lp_opamp_p_to_tempsense tempsense right_lp_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x33 vssa0 right_instramp_p_to_tempsense tempsense right_instramp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x1 vssa0 ulpcomp_p_to_tempsense tempsense ulpcomp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x3 vssa0 comp_p_to_tempsense tempsense comp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x5 vssa0 adc0_to_tempsense tempsense adc0 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x6 vssa0 ulpcomp_n_to_right_vref right_vref ulpcomp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x10 vssa0 comp_n_to_right_vref right_vref comp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x11 vssa0 adc1_to_right_vref right_vref adc1 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x12 vssa0 ulpcomp_p_to_left_vref left_vref ulpcomp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x14 vssa0 comp_p_to_left_vref left_vref comp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x16 vssa0 adc0_to_left_vref left_vref adc0 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x20 vssa0 ulpcomp_n_to_vinref vinref ulpcomp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x27 vssa0 comp_n_to_vinref vinref comp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x30 vssa0 adc1_to_vinref vinref adc1 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x32 vssa0 ulpcomp_p_to_voutref voutref ulpcomp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x34 vssa0 comp_p_to_voutref voutref comp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x35 vssa0 adc0_to_voutref voutref adc0 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x36 vssa0 right_instramp_p_to_left_vref left_vref right_instramp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x37 vssa0 right_hgbw_opamp_p_to_left_vref left_vref right_hgbw_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x38 vssa0 right_lp_opamp_p_to_left_vref left_vref right_lp_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x39 vssa0 left_lp_opamp_p_to_left_vref left_vref left_lp_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x40 vssa0 left_hgbw_opamp_p_to_left_vref left_vref left_hgbw_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x41 vssa0 left_instramp_p_to_left_vref left_vref left_instramp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x42 vssa0 right_instramp_n_to_vinref vinref right_instramp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x43 vssa0 right_hgbw_opamp_n_to_vinref vinref right_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x44 vssa0 right_lp_opamp_n_to_vinref vinref right_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x45 vssa0 left_lp_opamp_n_to_vinref vinref left_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x46 vssa0 left_hgbw_opamp_n_to_vinref vinref left_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x47 vssa0 left_instramp_n_to_vinref vinref left_instramp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x48 vssa0 right_instramp_p_to_voutref voutref right_instramp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x49 vssa0 right_hgbw_opamp_p_to_voutref voutref right_hgbw_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x50 vssa0 right_lp_opamp_p_to_voutref voutref right_lp_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x51 vssa0 left_lp_opamp_p_to_voutref voutref left_lp_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x52 vssa0 left_hgbw_opamp_p_to_voutref voutref left_hgbw_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x53 vssa0 left_instramp_p_to_voutref voutref left_instramp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
.ends


* expanding   symbol:  simple_switch_array_14.sym # of pins=34
** sym_path: /home/tim/gits/frigate_analog/xschem/simple_switch_array_14.sym
** sch_path: /home/tim/gits/frigate_analog/xschem/simple_switch_array_14.sch
.subckt simple_switch_array_14 vdda0 vssa0 vccd0 vssd0 right_hgbw_opamp_n_to_dac1 right_hgbw_opamp_p_to_dac0 right_hgbw_opamp_n
+ right_hgbw_opamp_p right_lp_opamp_n_to_dac1 right_lp_opamp_p_to_dac0 right_lp_opamp_n right_lp_opamp_p left_hgbw_opamp_n left_hgbw_opamp_p
+ left_lp_opamp_n_to_dac1 left_lp_opamp_p_to_dac0 left_lp_opamp_n left_lp_opamp_p ulpcomp_p ulpcomp_n left_hgbw_opamp_n_to_dac1 left_hgbw_opamp_p_to_dac0
+ comp_p comp_n adc0 adc1 ulpcomp_n_to_dac1 ulpcomp_p_to_dac0 dac0 dac1 comp_n_to_dac1 comp_p_to_dac0 adc1_to_dac1 adc0_to_dac0
*.PININFO vccd0:B vdda0:B vssa0:B vssd0:B right_hgbw_opamp_n_to_dac1:I right_lp_opamp_n_to_dac1:I left_lp_opamp_n_to_dac1:I
*+ left_hgbw_opamp_n_to_dac1:I ulpcomp_p_to_dac0:I comp_p_to_dac0:I adc0_to_dac0:I dac1:B right_hgbw_opamp_p_to_dac0:I right_lp_opamp_p_to_dac0:I
*+ left_lp_opamp_p_to_dac0:I left_hgbw_opamp_p_to_dac0:I ulpcomp_n_to_dac1:I comp_n_to_dac1:I adc1_to_dac1:I dac0:B right_hgbw_opamp_n:B right_hgbw_opamp_p:B
*+ right_lp_opamp_n:B right_lp_opamp_p:B left_hgbw_opamp_n:B left_hgbw_opamp_p:B left_lp_opamp_n:B left_lp_opamp_p:B ulpcomp_p:B ulpcomp_n:B comp_p:B
*+ comp_n:B adc0:B adc1:B
x2 vssa0 right_hgbw_opamp_n_to_dac1 dac1 right_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x3 vssa0 right_lp_opamp_n_to_dac1 dac1 right_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x4 vssa0 left_lp_opamp_n_to_dac1 dac1 left_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x5 vssa0 left_hgbw_opamp_n_to_dac1 dac1 left_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x7 vssa0 ulpcomp_p_to_dac0 dac0 ulpcomp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x8 vssa0 comp_p_to_dac0 dac0 comp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x9 vssa0 adc0_to_dac0 dac0 adc0 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x12 vssa0 right_hgbw_opamp_p_to_dac0 dac0 right_hgbw_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x13 vssa0 right_lp_opamp_p_to_dac0 dac0 right_lp_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x14 vssa0 left_lp_opamp_p_to_dac0 dac0 left_lp_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x15 vssa0 left_hgbw_opamp_p_to_dac0 dac0 left_hgbw_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x17 vssa0 ulpcomp_n_to_dac1 dac1 ulpcomp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x18 vssa0 comp_n_to_dac1 dac1 comp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x19 vssa0 adc1_to_dac1 dac1 adc1 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
.ends


* expanding   symbol:  simple_switch_array_16.sym # of pins=38
** sym_path: /home/tim/gits/frigate_analog/xschem/simple_switch_array_16.sym
** sch_path: /home/tim/gits/frigate_analog/xschem/simple_switch_array_16.sch
.subckt simple_switch_array_16 vdda0 vssa0 vccd0 vssd0 right_instramp_n_to_sio1 right_instramp_p_to_sio0 sio0 sio1
+ right_hgbw_opamp_n_to_sio1 right_hgbw_opamp_p_to_sio0 right_instramp_n right_instramp_p right_hgbw_opamp_n right_hgbw_opamp_p right_lp_opamp_n_to_sio1
+ right_lp_opamp_n right_lp_opamp_p_to_sio0 right_lp_opamp_p left_instramp_n left_instramp_p left_hgbw_opamp_n left_lp_opamp_n_to_sio1
+ left_lp_opamp_p_to_sio0 left_hgbw_opamp_p left_lp_opamp_n left_lp_opamp_p ulpcomp_p left_hgbw_opamp_n_to_sio1 left_hgbw_opamp_p_to_sio0 ulpcomp_n comp_p
+ comp_n left_instramp_n_to_sio1 left_instramp_p_to_sio0 ulpcomp_n_to_sio1 ulpcomp_p_to_sio0 comp_n_to_sio1 comp_p_to_sio0
*.PININFO vccd0:B vdda0:B vssa0:B vssd0:B right_hgbw_opamp_n_to_sio1:I right_lp_opamp_n_to_sio1:I left_lp_opamp_n_to_sio1:I
*+ left_hgbw_opamp_n_to_sio1:I ulpcomp_p_to_sio0:I comp_p_to_sio0:I sio1:B right_hgbw_opamp_p_to_sio0:I right_lp_opamp_p_to_sio0:I left_lp_opamp_p_to_sio0:I
*+ left_hgbw_opamp_p_to_sio0:I ulpcomp_n_to_sio1:I comp_n_to_sio1:I sio0:B right_hgbw_opamp_n:B right_hgbw_opamp_p:B right_lp_opamp_n:B right_lp_opamp_p:B
*+ left_hgbw_opamp_n:B left_hgbw_opamp_p:B left_lp_opamp_n:B left_lp_opamp_p:B ulpcomp_p:B ulpcomp_n:B comp_p:B comp_n:B right_instramp_n_to_sio1:I
*+ right_instramp_p_to_sio0:I left_instramp_n_to_sio1:I left_instramp_p_to_sio0:I right_instramp_n:B right_instramp_p:B left_instramp_n:B left_instramp_p:B
x2 vssa0 right_hgbw_opamp_n_to_sio1 sio1 right_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x3 vssa0 right_lp_opamp_n_to_sio1 sio1 right_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x4 vssa0 left_lp_opamp_n_to_sio1 sio1 left_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x5 vssa0 left_hgbw_opamp_n_to_sio1 sio1 left_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x7 vssa0 ulpcomp_p_to_sio0 sio0 ulpcomp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x8 vssa0 comp_p_to_sio0 sio0 comp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x12 vssa0 right_hgbw_opamp_p_to_sio0 sio0 right_hgbw_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x13 vssa0 right_lp_opamp_p_to_sio0 sio0 right_lp_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x14 vssa0 left_lp_opamp_p_to_sio0 sio0 left_lp_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x15 vssa0 left_hgbw_opamp_p_to_sio0 sio0 left_hgbw_opamp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x17 vssa0 ulpcomp_n_to_sio1 sio1 ulpcomp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x18 vssa0 comp_n_to_sio1 sio1 comp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x1 vssa0 right_instramp_n_to_sio1 sio1 right_instramp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x6 vssa0 right_instramp_p_to_sio0 sio0 right_instramp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x9 vssa0 left_instramp_n_to_sio1 sio1 left_instramp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x10 vssa0 left_instramp_p_to_sio0 sio0 left_instramp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
.ends


* expanding   symbol:  user_switch_array_15.sym # of pins=49
** sym_path: /home/tim/gits/frigate_analog/xschem/user_switch_array_15.sym
** sch_path: /home/tim/gits/frigate_analog/xschem/user_switch_array_15.sch
.subckt user_switch_array_15 user_to_comp_n[1] user_to_comp_n[0] user_to_comp_p[1] user_to_comp_p[0] vdda0 user_to_ulpcomp_n[1]
+ user_to_ulpcomp_n[0] vssa0 vccd0 user_to_ulpcomp_p[1] user_to_ulpcomp_p[0] vssd0 user_to_adc0[1] user_to_adc0[0] user_to_adc1[1] user_to_adc1[0]
+ vbgtc_to_user user_comp_n comp_n user_vbgtc vbgtc vbgsc_to_user user_comp_p comp_p user_vbgsc vbgsc dac0_to_user user_ulpcomp_n ulpcomp_n
+ user_dac0 dac0 dac1_to_user user_ulpcomp_p ulpcomp_p user_dac1 dac1 tempsense_to_user user_adc0 adc0 user_tempsense tempsense
+ right_vref_to_user user_adc1 adc1 user_right_vref right_vref left_vref_to_user user_left_vref left_vref vinref_to_user user_vinref vinref
+ voutref_to_user user_voutref voutref
*.PININFO vccd0:B vdda0:B vssa0:B vssd0:B vbgtc_to_user:I vbgsc_to_user:I dac0_to_user:I dac1_to_user:I vinref_to_user:I
*+ voutref_to_user:I tempsense_to_user:I right_vref_to_user:I left_vref_to_user:I ulpcomp_p:B ulpcomp_n:B comp_p:B comp_n:B adc0:B adc1:B dac0:B
*+ dac1:B tempsense:B right_vref:B left_vref:B vinref:B voutref:B vbgsc:B vbgtc:B user_vbgtc:B user_vbgsc:B user_dac0:B user_dac1:B
*+ user_tempsense:B user_right_vref:B user_left_vref:B user_vinref:B user_voutref:B user_adc1:B user_adc0:B user_ulpcomp_p:B user_ulpcomp_n:B
*+ user_comp_p:B user_comp_n:B user_to_comp_n[1:0]:I user_to_comp_p[1:0]:I user_to_ulpcomp_n[1:0]:I user_to_ulpcomp_p[1:0]:I user_to_adc0[1:0]:I
*+ user_to_adc1[1:0]:I
x2 vssa0 vbgtc_to_user user_vbgtc vbgtc vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x3 vssa0 vbgsc_to_user user_vbgsc vbgsc vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x4 vssa0 dac0_to_user user_dac0 dac0 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x5 vssa0 dac1_to_user user_dac1 dac1 vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x8 vssa0 vinref_to_user user_vinref vinref vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x9 vssa0 voutref_to_user user_voutref voutref vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x17 vssa0 tempsense_to_user user_tempsense tempsense vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x18 vssa0 right_vref_to_user user_right_vref right_vref vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x19 vssa0 left_vref_to_user user_left_vref left_vref vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x13 vssa0 user_to_adc1[0] user_adc1 adc1 vdda0 vccd0 vssd0 user_to_adc1[1] isolated_switch_large
x1 vssa0 user_to_adc0[0] user_adc0 adc0 vdda0 vccd0 vssd0 user_to_adc0[1] isolated_switch_large
x6 vssa0 user_to_ulpcomp_p[0] user_ulpcomp_p ulpcomp_p vdda0 vccd0 vssd0 user_to_ulpcomp_p[1] isolated_switch_large
x7 vssa0 user_to_ulpcomp_n[0] user_ulpcomp_n ulpcomp_n vdda0 vccd0 vssd0 user_to_ulpcomp_n[1] isolated_switch_large
x10 vssa0 user_to_comp_p[0] user_comp_p comp_p vdda0 vccd0 vssd0 user_to_comp_p[1] isolated_switch_large
x11 vssa0 user_to_comp_n[0] user_comp_n comp_n vdda0 vccd0 vssd0 user_to_comp_n[1] isolated_switch_large
.ends


* expanding   symbol:  simple_switch_array_12.sym # of pins=32
** sym_path: /home/tim/gits/frigate_analog/xschem/simple_switch_array_12.sym
** sch_path: /home/tim/gits/frigate_analog/xschem/simple_switch_array_12.sch
.subckt simple_switch_array_12 vdda0 vssa0 vccd0 vssd0 right_instramp_p_to_right_rheostat1_out
+ right_instramp_n_to_right_rheostat1_out right_rheostat1_in right_hgbw_opamp_n left_instramp_p_to_left_rheostat1_out right_hgbw_opamp_n_to_rheostat_tap right_lp_opamp_n
+ right_rheostat1_tap left_hgbw_opamp_n right_instramp_p_to_left_rheostat2_out left_instramp_n_to_left_rheostat1_out left_lp_opamp_n right_rheostat2_in
+ right_lp_opamp_n_to_rheostat_tap left_instramp_p_to_right_rheostat2_out right_rheostat2_tap right_instramp_n_to_left_rheostat2_out left_rheostat2_in
+ left_lp_opamp_n_to_rheostat_tap left_rheostat2_tap left_instramp_n_to_right_rheostat2_out left_rheostat1_in left_hgbw_opamp_n_to_rheostat_tap left_rheostat1_tap
+ left_instramp_n left_instramp_p right_instramp_n right_instramp_p
*.PININFO vccd0:B vdda0:B vssa0:B vssd0:B right_instramp_n_to_right_rheostat1_out:I left_instramp_n_to_right_rheostat2_out:I
*+ right_instramp_n_to_left_rheostat2_out:I left_instramp_n_to_left_rheostat1_out:I right_instramp_p_to_right_rheostat1_out:I left_instramp_p_to_right_rheostat2_out:I
*+ right_instramp_p_to_left_rheostat2_out:I left_instramp_p_to_left_rheostat1_out:I right_hgbw_opamp_n:B right_lp_opamp_n:B left_hgbw_opamp_n:B left_lp_opamp_n:B
*+ right_lp_opamp_n_to_rheostat_tap:I right_hgbw_opamp_n_to_rheostat_tap:I left_hgbw_opamp_n_to_rheostat_tap:I left_lp_opamp_n_to_rheostat_tap:I right_rheostat1_in:B
*+ right_rheostat1_tap:B right_rheostat2_in:B right_rheostat2_tap:B left_rheostat2_in:B left_rheostat2_tap:B left_rheostat1_in:B left_rheostat1_tap:B
*+ right_instramp_n:B right_instramp_p:B left_instramp_n:B left_instramp_p:B
x2 vssa0 right_instramp_n_to_right_rheostat1_out right_rheostat1_in right_instramp_n vdda0 vccd0 vssd0
+ simplest_analog_switch_ena1v8
x3 vssa0 left_instramp_n_to_right_rheostat2_out right_rheostat2_in left_instramp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x4 vssa0 right_instramp_n_to_left_rheostat2_out left_rheostat2_in right_instramp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x5 vssa0 left_instramp_n_to_left_rheostat1_out left_rheostat1_in left_instramp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x7 vssa0 left_lp_opamp_n_to_rheostat_tap left_rheostat2_tap left_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x8 vssa0 left_hgbw_opamp_n_to_rheostat_tap left_rheostat1_tap left_hgbw_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x12 vssa0 right_instramp_p_to_right_rheostat1_out right_rheostat1_in right_instramp_p vdda0 vccd0 vssd0
+ simplest_analog_switch_ena1v8
x13 vssa0 left_instramp_p_to_right_rheostat2_out right_rheostat2_in left_instramp_p vdda0 vccd0 vssd0
+ simplest_analog_switch_ena1v8
x14 vssa0 right_instramp_p_to_left_rheostat2_out left_rheostat2_in right_instramp_p vdda0 vccd0 vssd0
+ simplest_analog_switch_ena1v8
x15 vssa0 left_instramp_p_to_left_rheostat1_out left_rheostat1_in left_instramp_p vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
x17 vssa0 right_hgbw_opamp_n_to_rheostat_tap right_rheostat1_tap right_hgbw_opamp_n vdda0 vccd0 vssd0
+ simplest_analog_switch_ena1v8
x18 vssa0 right_lp_opamp_n_to_rheostat_tap right_rheostat2_tap right_lp_opamp_n vdda0 vccd0 vssd0 simplest_analog_switch_ena1v8
.ends


* expanding   symbol:  switch_array_2.sym # of pins=10
** sym_path: /home/tim/gits/frigate_analog/xschem/switch_array_2.sym
** sch_path: /home/tim/gits/frigate_analog/xschem/switch_array_2.sch
.subckt switch_array_2 avdd dvdd dvss avss channel0_out channel0_in_to_out[1] channel0_in_to_out[0] channel0_in
+ channel1_in_to_out[1] channel1_in_to_out[0] channel1_out channel1_in
*.PININFO channel0_in:B avdd:B dvdd:B dvss:B avss:B channel0_in_to_out[1:0]:I channel0_out:B channel1_in:B channel1_out:B
*+ channel1_in_to_out[1:0]:I
x1 avss channel0_in_to_out[0] channel0_out channel0_in avdd dvdd dvss channel0_in_to_out[1] isolated_switch_xlarge
x2 avss channel1_in_to_out[0] channel1_out channel1_in avdd dvdd dvss channel1_in_to_out[1] isolated_switch_xlarge
.ends


* expanding   symbol:  simple_analog_mux_sel1v8.sym # of pins=8
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_mux_sel1v8.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_mux_sel1v8.sch
.subckt simple_analog_mux_sel1v8 avss selA inA avdd inB out dvdd dvss
*.PININFO selA:I avss:B out:B inA:B avdd:B dvdd:B dvss:B inB:B
x2 selA dvdd dvss dvss avdd avdd net3 sky130_fd_sc_hvl__lsbuflv2hv_1
x3 net1 net2 avss out inA avdd simple_analog_switch_2
x1 net3 dvss dvss avdd avdd net2 sky130_fd_sc_hvl__inv_2
x4 net2 dvss dvss avdd avdd net1 sky130_fd_sc_hvl__inv_2
x5[1] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x5[0] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x5 net2 net1 avss inB out avdd simple_analog_switch_2
x6 selA dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
.ends


* expanding   symbol:  sky130_ef_ip__idac3v_8bit.sym # of pins=11
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/sky130_ef_ip__idac3v_8bit.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/sky130_ef_ip__idac3v_8bit.sch
.subckt sky130_ef_ip__idac3v_8bit ena ref_in vbg ref_sel_vbg dvdd dvss avdd din[7] din[6] din[5] din[4] din[3] din[2] din[1]
+ din[0] avss src_out snk_out
*.PININFO ena:I din[7:0]:I ref_sel_vbg:I vbg:I ref_in:I src_out:B snk_out:B dvdd:B dvss:B avdd:B avss:B
x1 avdd ena vbg net4 avss dvdd dvss ref_sel_vbg ref_in dvss net2 net1 net3 net5 dvss bias_generator_fe
x2 dvdd dvss din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] avdd net1 net3 src_out snk_out net2 avss
+ bias_generator_idac_be
* noconn #net4
* noconn #net5
.ends


* expanding   symbol:  sky130_ajc_ip__brownout.sym # of pins=22
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ajc_ip__brownout/xschem/sky130_ajc_ip__brownout.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ajc_ip__brownout/xschem/sky130_ajc_ip__brownout.sch
.subckt sky130_ajc_ip__brownout avdd avss outb dvdd osc_ck dvss dcomp vbg_1v2 otrip[2] otrip[1] otrip[0] itest brout_filt vtrip[2]
+ vtrip[1] vtrip[0] vin_brout ena force_ena_rc_osc vin_vunder force_dis_rc_osc timed_out vunder force_short_oneshot isrc_sel ibg_200n
*.PININFO avdd:I avss:I dvdd:I dvss:I vbg_1v2:I otrip[2:0]:I ena:I force_dis_rc_osc:I force_short_oneshot:I isrc_sel:I ibg_200n:I
*+ vin_brout:O outb:O osc_ck:O brout_filt:O itest:O timed_out:O vtrip[2:0]:I vin_vunder:O vunder:O force_ena_rc_osc:I dcomp:O
xIana vin_brout otrip_decoded_7_ otrip_decoded_6_ otrip_decoded_5_ otrip_decoded_4_ otrip_decoded_3_ otrip_decoded_2_
+ otrip_decoded_1_ otrip_decoded_0_ vin_vunder vbg_1v2 ena avdd ibg_200n itest avss dvdd isrc_sel dvss vtrip_decoded_7_ vtrip_decoded_6_
+ vtrip_decoded_5_ vtrip_decoded_4_ vtrip_decoded_3_ vtrip_decoded_2_ vtrip_decoded_1_ vtrip_decoded_0_ dcomp brout_filt osc_ck osc_ena vunder outb
+ outb_unbuf brownout_ana
xIdig brout_filt dcomp ena force_dis_rc_osc force_ena_rc_osc force_short_oneshot osc_ck osc_ena outb_unbuf timed_out dvdd dvss
+ otrip[2] otrip[1] otrip[0] otrip_decoded_7_ otrip_decoded_6_ otrip_decoded_5_ otrip_decoded_4_ otrip_decoded_3_ otrip_decoded_2_
+ otrip_decoded_1_ otrip_decoded_0_ vtrip[2] vtrip[1] vtrip[0] vtrip_decoded_7_ vtrip_decoded_6_ vtrip_decoded_5_ vtrip_decoded_4_ vtrip_decoded_3_
+ vtrip_decoded_2_ vtrip_decoded_1_ vtrip_decoded_0_ brownout_dig
XMdum0 otrip[2] dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XMdum1 otrip[1] dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XMdum2 otrip[0] dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XMdum3 vtrip[2] dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XMdum4 vtrip[1] dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XMdum5 vtrip[0] dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XMdum6 ena dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XMdum7 force_ena_rc_osc dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XMdum8 force_dis_rc_osc dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XMdum9 force_short_oneshot dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XMdum10 vbg_1v2 dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XMdum11 isrc_sel dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XMdum12 vin_brout dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
XMdum13 vin_vunder dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=2
.ends


* expanding   symbol:  sky130_iic_ip__audiodac_drv_lite.sym # of pins=7
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_iic_ip__audiodac_lite/xschem/sky130_iic_ip__audiodac_drv_lite.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_iic_ip__audiodac_lite/xschem/sky130_iic_ip__audiodac_drv_lite.sch
.subckt sky130_iic_ip__audiodac_drv_lite out_p vdd in_hi in_p in_n vss out_n
*.PININFO in_p:I in_n:I out_p:O out_n:O vdd:I in_hi:I vss:I
x1 vdd drv_p drv_n in_hi in_p in_n vss audiodac_drv_ls
x2 vdd net1 net2 vss audiodac_drv_latch
XMdecouple vdd vss vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=10 W=55 nf=1 m=2
x5 vdd drv_p out_p vss net1 audiodac_drv_lite_half
x6 vdd drv_n out_n vss net2 audiodac_drv_lite_half
.ends


* expanding   symbol:  sky130_pa_ip__instramp.sym # of pins=10
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/sky130_pa_ip__instramp.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/sky130_pa_ip__instramp.sch
.subckt sky130_pa_ip__instramp V[9] V[8] V[7] V[6] V[5] V[4] V[3] V[2] V[1] V[0] VCM IBIAS AVDD VINN DVDD VOUT AVSS DVSS VINP
*.PININFO VCM:I AVDD:B VOUT:O IBIAS:I DVDD:B AVSS:B DVSS:B V[9:0]:I VINP:I VINN:I
x1 V[6] V[5] V[8] V[9] V[7] VO1 DVDD AVDD VOUT V[4] V[3] V[2] V[1] V[0] VCM DVSS AVSS VBIAS Parallel_10B_Block2
x2 net1 VINP VO1 VINN VCM AVSS VBIAS Input_Stage_v1
VI2 AVDD net1 0
.save i(vi2)
x3 VBIAS IBIAS AVSS vbias_gen_pga
.ends


* expanding   symbol:  sky130_ef_ip__scomp3v.sym # of pins=8
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__ccomp3v/xschem/sky130_ef_ip__scomp3v.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__ccomp3v/xschem/sky130_ef_ip__scomp3v.sch
.subckt sky130_ef_ip__scomp3v VOUT DVDD DVSS VDD VSS VINP VINM ENA
*.PININFO VDD:I VOUT:O VSS:I VINP:I VINM:I DVDD:I DVSS:I ENA:I
x3 ENA DVDD DVSS DVSS VDD VDD ena3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x1 VDD VBN VSS VINP VOUT VINM DVDD ena3v3 DVSS comparator_high_gain
x2 VDD VSS VBN ena3v3 scomp_bias
x4 ENA DVSS DVSS VDD VDD sky130_fd_sc_hvl__diode_2
.ends


* expanding   symbol:  sky130_td_ip__opamp_hp_narrow.sym # of pins=9
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_td_ip__opamp_hp/xschem/sky130_td_ip__opamp_hp_narrow.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_td_ip__opamp_hp/xschem/sky130_td_ip__opamp_hp_narrow.sch
.subckt sky130_td_ip__opamp_hp_narrow avdd vout ibias vinn vinp avss dvdd dvss ena
*.PININFO vinn:I vinp:I vout:O ena:I ibias:I avss:I avdd:I dvdd:I dvss:I
XM3 net45 vinn vtailn avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=24
XM4 net46 vinp vtailn avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=24
XMB3 vtailn vb3 net12 avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=4.5 nf=1 m=16
XMB4 net12 vb4 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=4.5 nf=1 m=16
XM1 net43 vinn vtailp avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=6 nf=1 m=24
XM2 net44 vinp vtailp avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=6 nf=1 m=24
XMB2 vtailp vb2 net11 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=9 nf=1 m=16
XMB1 net11 vb1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=9 nf=1 m=16
XM12 net4 net5 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=12 nf=1 m=18
XM11 net3 net5 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=12 nf=1 m=18
XM14 net7 vb2 net4 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=12 nf=1 m=18
XM13 net5 vb2 net3 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=12 nf=1 m=18
XM18 net2 net6 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=6 nf=1 m=12
XM16 net55 vb3 net2 avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=6 nf=1 m=12
XM17 net1 net6 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=6 nf=1 m=12
XM15 net6 vb3 net1 avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=6 nf=1 m=12
XM28 net19 net9 net5 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=4.2 nf=1 m=6
XM27 net5 net10 net19 avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=2 nf=1 m=6
XM20 net8 net9 net7 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4.2 nf=2 m=3
XM19 net7 net10 net8 avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=2 nf=1 m=3
XM26 vout net8 net36 net36 sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=10 nf=1 m=32
XM25 vout net7 net37 net37 sky130_fd_pr__pfet_g5v0d10v5 L=1 W=25 nf=1 m=32
XMB9 ibias net33 net34 avss sky130_fd_pr__nfet_g5v0d10v5 L=2.0 W=2 nf=1 m=2
XMB11 net34 net31 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2.0 W=2 nf=1 m=2
XMB10 net53 net33 net20 avss sky130_fd_pr__nfet_g5v0d10v5 L=2.0 W=2 nf=1 m=10
XMB12 net20 net31 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2.0 W=2 nf=1 m=10
XMB15 net21 net38 net32 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=2 nf=1 m=2
XMB13 net32 net22 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=2 nf=1 m=2
XMB16 net39 net38 net23 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=2 nf=1 m=8
XMB14 net23 net22 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=2 nf=1 m=8
XMB17 vb7 vb7 vb8 avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=2 nf=1 m=2
XMB19 vb8 vb8 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=2 nf=1 m=2
XMB18 net50 vb7 net24 avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=2 nf=1 m=10
XMB20 net24 vb8 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=2 nf=1 m=10
XMB22 net51 vb7 net25 avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=2 nf=1 m=10
XMB23 net25 vb8 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=2 nf=1 m=10
XMB21 vb2 vb2 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=3 nf=1 m=1
XMB27 vb6 vb6 vb5 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=4 nf=1 m=6
XMB24 vb5 vb5 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=4 nf=1 m=6
XMB28 net40 vb6 net26 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=4 nf=1 m=6
XMB25 net26 vb5 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=4 nf=1 m=6
XMB29 net41 vb6 net27 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=4 nf=1 m=12
XMB26 net27 vb5 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=4 nf=1 m=12
XMB30 vb3 vb3 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=1.5 nf=1 m=1
XMB31 vb4 vb3 net28 avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=4.5 nf=1 m=4
XMB33 net28 vb4 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=4.5 nf=1 m=4
XMB32 net52 vb3 net29 avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=4.5 nf=1 m=4
XMB34 net29 vb4 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=4.5 nf=1 m=4
XM36 vb1 vb2 net30 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=9 nf=1 m=4
XMB35 net30 vb1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=9 nf=1 m=4
XM24 net14 net14 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=2 nf=1 m=4
XM23 net10 net10 net14 avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=2 nf=1 m=4
XMB5 net13 vb5 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=4 nf=1 m=6
XMB6 net10 vb6 net13 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=4 nf=1 m=6
XM21 net15 net15 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=4 nf=1 m=4
XM22 net9 net9 net15 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1.0 W=4 nf=1 m=4
XMB8 net16 vb8 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=2 nf=1 m=10
XMB7 net9 vb7 net16 avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=2 nf=1 m=10
XM5 net54 vb3 vtailn avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4.5 nf=1 m=8
XM6 net18 net18 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=16 nf=1 m=4
XM7 vtailp net18 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=16 nf=1 m=12
XM8 net42 vb2 vtailp avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=9 nf=1 m=8
XM9 net17 net17 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=8 nf=1 m=4
XM10 vtailn net17 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=8 nf=1 m=12
V_ID1 net43 net1 0
.save i(v_id1)
V_ID2 net44 net2 0
.save i(v_id2)
V_ID3 net3 net45 0
.save i(v_id3)
V_ID4 net4 net46 0
.save i(v_id4)
V_ID25 avdd net37 0
.save i(v_id25)
V_ID26 net36 avss 0
.save i(v_id26)
XM29 net47 net35 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=4
XM30 net35 net47 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=4
XM31 net47 net48 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=2
XM32 net35 net49 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=2
XM33 net49 net48 dvss dvss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM34 net49 net48 dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM35 net11 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM40 net12 enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM41 net1 enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM37 net16 enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM38 net17 enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM42 net13 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM43 net18 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM44 net34 ena_avdd net31 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM45 net20 enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM50 net23 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM54 net48 ena dvss dvss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM55 net48 ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM56 ena_avdd net35 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM57 ena_avdd net35 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM58 enab_avdd net47 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM59 enab_avdd net47 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM60 vb1 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM61 net5 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM62 vb4 enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM63 net6 enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM64 net2 enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM65 net3 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM66 net4 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM67 net31 enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM68 net22 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM69 vb8 enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM70 vb5 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM71 vb7 enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM72 vb6 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM73 net10 enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM74 net9 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM75 vb2 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM76 vb3 enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
V_IB1 net21 net53 0
.save i(v_ib1)
V_IB2 net39 vb7 0
.save i(v_ib2)
V_IB3 vb2 net50 0
.save i(v_ib3)
V_IB4 vb6 net51 0
.save i(v_ib4)
V_IB5 net40 vb3 0
.save i(v_ib5)
V_IB6 net41 vb4 0
.save i(v_ib6)
V_IB7 vb1 net52 0
.save i(v_ib7)
XM78 net32 enab_avdd net22 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM79 net32 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM81 net21 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
V_ID9 net42 net17 0
.save i(v_id9)
V_ID6 net18 net54 0
.save i(v_id6)
V_ID15 net19 net6 0
.save i(v_id15)
V_ID16 net8 net55 0
.save i(v_id16)
XM77 net7 ena_avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM82 vinn enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM83 vinp enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM80 ibias ena_avdd net33 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM84 net21 enab_avdd net38 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM85 net33 enab_avdd avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XC3 net8 resb_in sky130_fd_pr__cap_mim_m3_1 W=12 L=12 m=9
XC1 net7 resa_in sky130_fd_pr__cap_mim_m3_1 W=12 L=12 m=9
XMB36 net20 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2.0 W=2 nf=1 m=2
XMB37 net34 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2.0 W=2 nf=1 m=2
XMB38 net20 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2.0 W=2 nf=1 m=2
XMB39 vtailn avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1.0 W=8 nf=1 m=2
XMB40 net35 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=2
XMB41 net18 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4.5 nf=1 m=2
XMB42 net12 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4.5 nf=1 m=2
XMB43 vb4 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4.5 nf=1 m=2
XMB44 vb1 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4.5 nf=1 m=2
XMB45 vtailn avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4.5 nf=1 m=2
XMB46 vtailn avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=4
XMB47 net6 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XMB48 net8 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XMB49 net7 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XMB50 net10 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XMB51 avss avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XMB52 net6 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=6 nf=1 m=2
XMB53 net8 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=6 nf=1 m=2
XMB54 avss avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=6 nf=1 m=2
XMB55 net25 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XMB56 net24 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XMB57 net16 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XMB58 vb7 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XMB59 net24 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XMB60 net25 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XMB61 net16 avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM39 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=2
XM46 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=16 nf=1 m=2
XM47 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=9 nf=1 m=2
XM48 vb1 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=9 nf=1 m=2
XM49 vtailp avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=9 nf=1 m=2
XM51 vtailp avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=6 nf=1 m=4
XM52 net5 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4.2 nf=1 m=2
XM53 net7 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4.2 nf=1 m=1
XM86 net8 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4.2 nf=1 m=1
XM87 net15 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM88 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM89 net5 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=12 nf=1 m=2
XM90 net7 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=12 nf=1 m=2
XM91 net4 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=12 nf=1 m=2
XM92 net32 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM93 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=2
XM94 vb7 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM95 net15 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM96 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=2
XM97 net26 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=2
XM98 net13 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=2
XM99 vb3 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=2
XM100 vb4 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=2
XM101 net10 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=2
XM102 vb6 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=2
XM103 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=25 nf=1 m=2
XR3 net56 resa_in avss sky130_fd_pr__res_high_po_0p69 L=1.4 mult=1 m=1
XR5 net56 vout avss sky130_fd_pr__res_high_po_0p69 L=1.4 mult=1 m=1
XR6 net57 resb_in avss sky130_fd_pr__res_high_po_0p69 L=1.4 mult=1 m=1
XR7 net57 vout avss sky130_fd_pr__res_high_po_0p69 L=1.4 mult=1 m=1
XR1 avss avss avss sky130_fd_pr__res_high_po_0p69 L=1.4 mult=1 m=1
XR2 avss avss avss sky130_fd_pr__res_high_po_0p69 L=1.4 mult=1 m=1
XMB62 avss avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=1 m=2
XM104 vtailp avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=9 nf=1 m=2
XD1 dvss ena sky130_fd_pr__diode_pw2nd_05v5 area=211.6e9 perim=1.84e6
XC2 resb_in net8 sky130_fd_pr__cap_mim_m3_2 W=12 L=12 m=9
XC4 resa_in net7 sky130_fd_pr__cap_mim_m3_2 W=12 L=12 m=9
.ends


* expanding   symbol:  sky130_cw_ip__bandgap_nobias.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_cw_ip/xschem/sky130_cw_ip__bandgap_nobias.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_cw_ip/xschem/sky130_cw_ip__bandgap_nobias.sch
.subckt sky130_cw_ip__bandgap_nobias vdd vbg vss bias trim[15] trim[14] trim[13] trim[12] trim[11] trim[10] trim[9] trim[8]
+ trim[7] trim[6] trim[5] trim[4] trim[3] trim[2] trim[1] trim[0] vsub
*.PININFO vsub:B vss:B vdd:B vbg:O trim[15:0]:I bias:B
x1 vdd vbg vss bias trim[15] trim[14] trim[13] trim[12] trim[11] trim[10] trim[9] trim[8] trim[7] trim[6] trim[5] trim[4] trim[3]
+ trim[2] trim[1] trim[0] bandgap
.ends


* expanding   symbol:  sky130_ef_ip__biasgen4.sym # of pins=52
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/sky130_ef_ip__biasgen4.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/sky130_ef_ip__biasgen4.sch
.subckt sky130_ef_ip__biasgen4 ena avdd avss ref_in dvdd vbg ref_sel_vbg dvss lp1_src_100 en_lp1_bias en_lp1_trim_p en_lp2_bias
+ lp2_src_100 en_lp2_trim_p en_hgbw1_bias hgbw1_src_100 en_hgbw1_trim_p hgbw2_src_100 en_hgbw2_bias en_hgbw2_trim_p instr1_src_100
+ en_instr1_bias en_instr1_trim_p instr2_src_100 en_instr2_bias en_instr2_trim_p lsxo_src_50 en_lsxo_bias hsxo_src_100 en_hsxo_bias en_hsxo_trim_p
+ en_hsxo_trim_n comp_src_400 en_comp_bias en_comp_trim_p en_comp_trim_n ov_src_600 en_ov_bias en_idac_bias idac_src_1000 en_brnout_bias
+ brnout_src_200 en_user1_bias user_src_50 en_user2_bias user_src_150 en_user2_trim_p en_user2_trim_n en_src_test test_src_500 en_snk_test
+ bandgap_snk_250
*.PININFO avdd:B avss:B dvdd:B dvss:B lp1_src_100:B lp2_src_100:B hgbw1_src_100:B hgbw2_src_100:B instr1_src_100:B
*+ instr2_src_100:B lsxo_src_50:B hsxo_src_100:B comp_src_400:B ov_src_600:B idac_src_1000:B brnout_src_200:B user_src_50:B user_src_150:B
*+ test_src_500:B ena:I ref_in:I vbg:I ref_sel_vbg:I en_lp1_bias:I en_lp1_trim_p:I en_lp2_bias:I en_lp2_trim_p:I en_hgbw1_bias:I en_hgbw1_trim_p:I
*+ en_hgbw2_bias:I en_hgbw2_trim_p:I en_instr1_bias:I en_instr2_bias:I en_instr1_trim_p:I en_instr2_trim_p:I en_lsxo_bias:I en_hsxo_bias:I
*+ en_hsxo_trim_p:I en_hsxo_trim_n:I en_comp_bias:I en_comp_trim_p:I en_comp_trim_n:I en_ov_bias:I en_idac_bias:I en_brnout_bias:I en_user1_bias:I
*+ en_user2_bias:I en_user2_trim_p:I en_user2_trim_n:I en_src_test:I en_snk_test:I bandgap_snk_250:B
x1 avdd ena vbg net1 avss dvdd dvss ref_sel_vbg ref_in dvss net5 net4 net3 net2 dvss bias_generator_fe
* noconn #net1
* noconn #net2
x3 dvdd dvss en_hsxo_bias en_comp_trim_n en_ov_bias avdd en_comp_bias net4 en_hsxo_trim_n net3 en_lp1_bias en_user2_trim_n
+ en_lp2_bias en_hgbw1_bias lp1_src_100 test_src_500 lp2_src_100 en_hgbw2_bias user_src_50 idac_src_1000 lsxo_src_50 hsxo_src_100 comp_src_400
+ hgbw2_src_100 ov_src_600 user_src_150 instr1_src_100 instr2_src_100 hgbw1_src_100 en_instr1_bias en_instr2_bias en_src_test en_lsxo_bias
+ en_snk_test net5 en_user1_bias avss en_idac_bias en_user2_bias en_comp_trim_p en_hsxo_trim_p en_user2_trim_p en_lp1_trim_p en_lp2_trim_p
+ en_hgbw1_trim_p en_hgbw2_trim_p en_instr1_trim_p en_instr2_trim_p brnout_src_200 en_brnout_bias bandgap_snk_250 bias_generator_be4
.ends


* expanding   symbol:  sky130_sw_ip__por.sym # of pins=7
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_sw_ip__por/xschem/sky130_sw_ip__por.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_sw_ip__por/xschem/sky130_sw_ip__por.sch
.subckt sky130_sw_ip__por por avss avdd dvdd porb dvss porb_h[1] porb_h[0]
*.PININFO avdd:B por:O avss:B dvdd:B porb:O porb_h[1:0]:O dvss:B
x1 Vinn Vinp RST avss net1 dvdd vo net6 comparator_final
XR1 avss Vinn avss sky130_fd_pr__res_xhigh_po_0p35 L=1000 mult=1 m=1
XR10 Vinn Vinp avss sky130_fd_pr__res_xhigh_po_0p35 L=72 mult=1 m=1
XR12 Vinp net3 avss sky130_fd_pr__res_xhigh_po_0p35 L=600 mult=1 m=1
x2 RST por dvdd dvss net2 porb porb_h[1] porb_h[0] net6 delayPulse_final
XM2 avdd avdd net4 avss sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 m=1
Vrbranch Vproc net3 0
.save i(vrbranch)
Vcomp avdd net1 0
.save i(vcomp)
Vpulse avdd net2 0
.save i(vpulse)
XM1 net4 avdd Vproc avss sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 m=1
XR2 net5 Vinp avss sky130_fd_pr__res_xhigh_po_0p35 L=72 mult=1 m=1
XM3 net5 vo Vinn avss sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 m=1
.ends


* expanding   symbol:  sbvfcm.sym # of pins=5
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ak_ip__cmos_vref/xschem/sbvfcm.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ak_ip__cmos_vref/xschem/sbvfcm.sch
.subckt sbvfcm vdd pbias nbias vx vss
*.PININFO vss:B vdd:B vx:B pbias:B nbias:B
XM3 net1 vbias_st vx vss sky130_fd_pr__nfet_01v8 L=2 W=100 nf=8 m=1
XM4 net2 vbias_st vss vss sky130_fd_pr__nfet_01v8 L=2 W=5 nf=1 m=1
XM5 pbias nbias net1 vss sky130_fd_pr__nfet_01v8 L=10 W=10 nf=1 m=1
XM6 vbias_st nbias net2 vss sky130_fd_pr__nfet_01v8 L=10 W=10 nf=1 m=1
XM7 pbias pbias net6 vdd sky130_fd_pr__pfet_01v8 L=10 W=5 nf=1 m=1
XM8 vbias_st pbias net7 vdd sky130_fd_pr__pfet_01v8 L=10 W=5 nf=1 m=1
XM10 net4 net3 vss vss sky130_fd_pr__nfet_01v8 L=10 W=5 nf=1 m=1
XM11 net3 vbias_st vss vss sky130_fd_pr__nfet_01v8 L=5 W=10 nf=1 m=1
XC1 net5 net3 sky130_fd_pr__cap_mim_m3_1 W=5 L=5 m=2
Vm_st1 pbias net4 0
.save i(vm_st1)
Vm_st2 vdd net5 0
.save i(vm_st2)
Vm_b1 vdd net6 0
.save i(vm_b1)
Vm_b2 vdd net7 0
.save i(vm_b2)
.ends


* expanding   symbol:  output_amp.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ak_ip__cmos_vref/xschem/output_amp.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ak_ip__cmos_vref/xschem/output_amp.sch
.subckt output_amp vdd vo vp vn ibias vss
*.PININFO vp:I vn:I ibias:I vo:O vss:I vdd:I
XM1 ibias ibias vss vss sky130_fd_pr__nfet_01v8 L=1 W=2.5 nf=1 m=1
XM2 net2 ibias vss vss sky130_fd_pr__nfet_01v8 L=1 W=5 nf=1 m=1
XM7 vo_pre net1 net4 vdd sky130_fd_pr__pfet_01v8 L=10 W=5 nf=1 m=1
XM4 net7 vn vcm vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=2 m=1
XM5 net8 vp vcm vss sky130_fd_pr__nfet_01v8 L=2 W=10 nf=2 m=1
XM6 net1 net1 net3 vdd sky130_fd_pr__pfet_01v8 L=10 W=5 nf=1 m=1
Vm_b1 vdd net3 0
.save i(vm_b1)
XM3 net6 ibias vss vss sky130_fd_pr__nfet_01v8 L=1 W=8 nf=1 m=1
XM8 vo vo_pre net5 vdd sky130_fd_pr__pfet_01v8 L=5 W=40 nf=2 m=1
Vm_op vdd net5 0
.save i(vm_op)
Vm_cm vcm net2 0
.save i(vm_cm)
Vm_b2 vdd net4 0
.save i(vm_b2)
XC2 vo vo_pre sky130_fd_pr__cap_mim_m3_1 W=5 L=5 m=10
Vm_on vo net6 0
.save i(vm_on)
XM9 net1 vn net7 vss sky130_fd_pr__nfet_05v0_nvt L=2 W=20 nf=2 m=1
XM10 vo_pre vp net8 vss sky130_fd_pr__nfet_05v0_nvt L=2 W=20 nf=2 m=1
.ends


* expanding   symbol:  trim_res.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ak_ip__cmos_vref/xschem/trim_res.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ak_ip__cmos_vref/xschem/trim_res.sch
.subckt trim_res A trim0 trim2 trim3 trim1 B
*.PININFO trim0:I trim1:I trim2:I trim3:I B:B A:B
XM1 A trim3 net3 B sky130_fd_pr__nfet_01v8 L=2 W=10 nf=1 m=1
XM2 net3 trim2 net2 B sky130_fd_pr__nfet_01v8 L=2 W=10 nf=1 m=1
XM3 net2 trim1 net1 B sky130_fd_pr__nfet_01v8 L=2 W=10 nf=1 m=1
XM4 net1 trim0 B B sky130_fd_pr__nfet_01v8 L=2 W=10 nf=1 m=1
XR1 B net1 B sky130_fd_pr__res_xhigh_po_0p69 L=3.45 mult=1 m=1
XR2 net1 net2 B sky130_fd_pr__res_xhigh_po_0p69 L=6.9 mult=1 m=1
XR3 net2 net3 B sky130_fd_pr__res_xhigh_po_0p69 L=13.8 mult=1 m=1
XR4 net3 A B sky130_fd_pr__res_xhigh_po_0p69 L=27.6 mult=1 m=1
.ends


* expanding   symbol:  level_shifter_up.sym # of pins=7
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ak_ip__comparator/xschem/level_shifter_up.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ak_ip__comparator/xschem/level_shifter_up.sch
.subckt level_shifter_up VDD_HV xb_hv x_hv x_lv GND_HV VDD_LV GND_LV
*.PININFO VDD_HV:I GND_HV:I x_lv:I x_hv:O xb_hv:O VDD_LV:I GND_LV:I
XM65 xb_hv x_lv GND_HV GND_HV sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM66 x_hv xb_lv GND_HV GND_HV sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM67 xb_hv x_hv VDD_HV VDD_HV sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=1
XM68 x_hv xb_hv VDD_HV VDD_HV sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=1
XM1 xb_lv x_lv GND_LV GND_LV sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM3 xb_lv x_lv VDD_LV VDD_LV sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
.ends


* expanding   symbol:  EF_BANK_CAP_12.sym # of pins=16
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_BANK_CAP_12.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_BANK_CAP_12.sch
.subckt EF_BANK_CAP_12 D8 D0 D4 VP1 D9 D5 D1 VP2 D2 D6 VSS D7 D3 D10 D11 Vref
*.PININFO D0:B D1:B D2:B D3:B D4:B D5:B D6:B D7:B D8:B D9:B VSS:B VP1:B VP2:B D10:B D11:B Vref:B
x4 VP1 VSS D0 D1 D2 D3 D4 D5 Vref EF_LSB_CAP
x1 D8 D10 D9 VP2 D6 VSS D7 D11 EF_MSB_CAP
x2 VP1 VP2 VSS EF_SC_CAP
.ends


* expanding   symbol:  EF_AMUX0201_ARRAY1.sym # of pins=31
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_AMUX0201_ARRAY1.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_AMUX0201_ARRAY1.sch
.subckt EF_AMUX0201_ARRAY1 D0 SELD0 D1 SELD1 SELD2 D2 SELD3 SELD4 D3 SELD5 D4 SELD6 SELD7 D5 SELD8 D6 SELD9 D7 D8 D9 VDD DVSS VH
+ VL VSS D10 D11 SELD10 SELD11 VCM RST
*.PININFO VDD:B DVSS:B VH:B VL:B SELD0:I SELD1:I SELD2:I SELD3:I SELD4:I SELD5:I SELD6:I SELD7:I SELD8:I SELD9:I VSS:B D0:B D1:B
*+ D2:B D3:B D4:B D5:B D6:B D7:B D8:B D9:B SELD10:I SELD11:I D10:B D11:B VCM:B RST:B
x2 VDD D0 VSS VH VL SELD0 DVSS VCM RST EF_AMUX21x
x1 VDD D1 VSS VH VL SELD1 DVSS VCM RST EF_AMUX21x
x3 VDD D2 VSS VH VL SELD2 DVSS VCM RST EF_AMUX21x
x4 VDD D3 VSS VH VL SELD3 DVSS VCM RST EF_AMUX21x
x5 VDD D4 VSS VH VL SELD4 DVSS VCM RST EF_AMUX21x
x8 VDD D5 VSS VH VL SELD5 DVSS VCM RST EF_AMUX21x
x9 VDD D6 VSS VH VL SELD6 DVSS VCM RST EF_AMUX21x
x10 VDD D7 VSS VH VL SELD7 DVSS VCM RST EF_AMUX21x
x11 VDD D8 VSS VH VL SELD8 DVSS VCM RST EF_AMUX21x
x12 VDD D9 VSS VH VL SELD9 DVSS VCM RST EF_AMUX21x
x6 VDD D10 VSS VH VL SELD10 DVSS VCM RST EF_AMUX21x
x7 VDD D11 VSS VH VL SELD11 DVSS VCM RST EF_AMUX21x
.ends


* expanding   symbol:  EF_SW_RST.sym # of pins=8
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_SW_RST.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_SW_RST.sch
.subckt EF_SW_RST VP1 VP2 AVDD AVSS HOLD VIN DVSS HOLDB
*.PININFO HOLD:I AVDD:B AVSS:B VP2:B VP1:B VIN:B DVSS:B HOLDB:I
x4 HOLDB HOLD AVSS VIN VP1 AVDD simple_analog_switch
x5 HOLDB HOLD AVSS VP2 VIN AVDD simple_analog_switch
.ends


* expanding   symbol:  cdac_lvlshift_array.sym # of pins=32
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/cdac_lvlshift_array.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/cdac_lvlshift_array.sch
.subckt cdac_lvlshift_array sel3 sel3_3p3 sel7_3p3 sel7 sel11_3p3 sel11 sel6 sel6_3p3 sel10 sel2_3p3 sel10_3p3 sel2 sel1_3p3
+ sel5_3p3 sel5 sel1 sel9 sel9_3p3 vdd3p3 vss sel0_3p3 sel4 sel4_3p3 sel8_3p3 sel8 vdd1p8 sel0 hold_3p3 hold rst_3p3 rst holdb_3p3
*.PININFO sel0:I vdd3p3:B vss:B vdd1p8:B rst:I sel0_3p3:O rst_3p3:O sel1:I sel1_3p3:O sel2:I sel2_3p3:O sel3:I sel3_3p3:O sel4:I
*+ sel4_3p3:O sel5:I sel5_3p3:O sel6:I sel6_3p3:O sel7:I sel7_3p3:O sel8:I sel8_3p3:O sel9:I sel9_3p3:O sel10:I sel10_3p3:O sel11:I sel11_3p3:O
*+ hold:I hold_3p3:O holdb_3p3:O
x19 rst vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__diode_2
x20 sel0 vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__diode_2
x1 sel1 vdd1p8 vss vss vdd3p3 vdd3p3 sel1_3p3 sky130_fd_sc_hvl__lsbuflv2hv_1
x2 sel1 vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__diode_2
x3 sel0 vdd1p8 vss vss vdd3p3 vdd3p3 sel0_3p3 sky130_fd_sc_hvl__lsbuflv2hv_1
x4 rst vdd1p8 vss vss vdd3p3 vdd3p3 rst_3p3 sky130_fd_sc_hvl__lsbuflv2hv_1
x5 sel2 vdd1p8 vss vss vdd3p3 vdd3p3 sel2_3p3 sky130_fd_sc_hvl__lsbuflv2hv_1
x6 sel2 vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__diode_2
x7 sel3 vdd1p8 vss vss vdd3p3 vdd3p3 sel3_3p3 sky130_fd_sc_hvl__lsbuflv2hv_1
x8 sel3 vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__diode_2
x9 sel4 vdd1p8 vss vss vdd3p3 vdd3p3 sel4_3p3 sky130_fd_sc_hvl__lsbuflv2hv_1
x10 sel4 vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__diode_2
x11 sel5 vdd1p8 vss vss vdd3p3 vdd3p3 sel5_3p3 sky130_fd_sc_hvl__lsbuflv2hv_1
x12 sel5 vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__diode_2
x13 sel6 vdd1p8 vss vss vdd3p3 vdd3p3 sel6_3p3 sky130_fd_sc_hvl__lsbuflv2hv_1
x14 sel6 vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__diode_2
x15 sel7 vdd1p8 vss vss vdd3p3 vdd3p3 sel7_3p3 sky130_fd_sc_hvl__lsbuflv2hv_1
x16 sel7 vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__diode_2
x17 sel8 vdd1p8 vss vss vdd3p3 vdd3p3 sel8_3p3 sky130_fd_sc_hvl__lsbuflv2hv_1
x18 sel8 vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__diode_2
x21 sel9 vdd1p8 vss vss vdd3p3 vdd3p3 sel9_3p3 sky130_fd_sc_hvl__lsbuflv2hv_1
x22 sel9 vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__diode_2
x23 sel10 vdd1p8 vss vss vdd3p3 vdd3p3 sel10_3p3 sky130_fd_sc_hvl__lsbuflv2hv_1
x24 sel10 vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__diode_2
x25 sel11 vdd1p8 vss vss vdd3p3 vdd3p3 sel11_3p3 sky130_fd_sc_hvl__lsbuflv2hv_1
x26 sel11 vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__diode_2
x27 hold vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__diode_2
x28 hold vdd1p8 vss vss vdd3p3 vdd3p3 hold_3p3 sky130_fd_sc_hvl__lsbuflv2hv_1
x29[14] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29[13] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29[12] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29[11] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29[10] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29[9] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29[8] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29[7] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29[6] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29[5] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29[4] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29[3] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29[2] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29[1] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29[0] vss vss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_4
x29 hold_3p3 vss vss vdd3p3 vdd3p3 holdb_3p3 sky130_fd_sc_hvl__inv_2
* noconn vdd3p3
* noconn vss
* noconn vdd1p8
.ends


* expanding   symbol:  rheo_half.sym # of pins=21
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rheostat_8bit/xschem/rheo_half.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rheostat_8bit/xschem/rheo_half.sch
.subckt rheo_half vdd vss b3 b4 b3b b4b b5 res_in b6 b0 dum_in b6b b5b b0b b1 b1b b2 b2b out res_out dum_out
*.PININFO res_in:B res_out:B out:B vdd:B vss:B b3:I b3b:I b5:I b5b:I b6:I b6b:I dum_out:B dum_in:B b4:I b4b:I b0:I b0b:I b1:I
*+ b1b:I b2:I b2b:I
x1 b2 b2b b1 b1b b0 b0b vdd net9 net8 net44 net16 vss net15 rheo_column
x2 b2 b2b b1 b1b b0 b0b vdd net10 net7 net43 net8 vss net9 rheo_column
x3 b2 b2b b1 b1b b0 b0b vdd net11 net6 net42 net7 vss net10 rheo_column
x4 b2 b2b b1 b1b b0 b0b vdd net12 net5 net41 net6 vss net11 rheo_column
x5 b2 b2b b1 b1b b0 b0b vdd net13 net4 net40 net5 vss net12 rheo_column
x6 b2 b2b b1 b1b b0 b0b vdd net14 net3 net39 net4 vss net13 rheo_column
x7 b2 b2b b1 b1b b0 b0b vdd net2 net1 net38 net3 vss net14 rheo_column
x8 b2 b2b b1 b1b b0 b0b vdd dum_in res_in net37 net1 vss net2 rheo_column
x9 b2 b2b b1 b1b b0 b0b vdd net25 net24 net52 res_out vss dum_out rheo_column
x10 b2 b2b b1 b1b b0 b0b vdd net26 net23 net51 net24 vss net25 rheo_column
x11 b2 b2b b1 b1b b0 b0b vdd net27 net22 net50 net23 vss net26 rheo_column
x12 b2 b2b b1 b1b b0 b0b vdd net28 net21 net49 net22 vss net27 rheo_column
x13 b2 b2b b1 b1b b0 b0b vdd net29 net20 net48 net21 vss net28 rheo_column
x14 b2 b2b b1 b1b b0 b0b vdd net30 net19 net47 net20 vss net29 rheo_column
x15 b2 b2b b1 b1b b0 b0b vdd net18 net17 net46 net19 vss net30 rheo_column
x16 b2 b2b b1 b1b b0 b0b vdd net15 net16 net45 net17 vss net18 rheo_column
x17 vdd b4 net31 net54 b4b vss passtrans
x18 vdd b4b net31 net53 b4 vss passtrans
x19 vdd b4 net32 net55 b4b vss passtrans
x20 vdd b4b net32 net56 b4 vss passtrans
x21 vdd b4 net33 net57 b4b vss passtrans
x22 vdd b4b net33 net58 b4 vss passtrans
x23 vdd b4 net34 net59 b4b vss passtrans
x24 vdd b4b net34 net60 b4 vss passtrans
x25 vdd b5b net36 net34 b5 vss passtrans
x26 vdd b5 net36 net33 b5b vss passtrans
x27 vdd b5b net35 net32 b5 vss passtrans
x28 vdd b5 net35 net31 b5b vss passtrans
x29 vdd b6b out net36 b6 vss passtrans
x30 vdd b6 out net35 b6b vss passtrans
x33 vdd b3b net60 net37 b3 vss passtrans
x31 vdd b3 net60 net38 b3b vss passtrans
x32 vdd b3b net59 net39 b3 vss passtrans
x34 vdd b3 net59 net40 b3b vss passtrans
x35 vdd b3b net58 net41 b3 vss passtrans
x36 vdd b3 net58 net42 b3b vss passtrans
x37 vdd b3b net57 net43 b3 vss passtrans
x38 vdd b3 net57 net44 b3b vss passtrans
x39 vdd b3b net56 net45 b3 vss passtrans
x40 vdd b3 net56 net46 b3b vss passtrans
x41 vdd b3b net55 net47 b3 vss passtrans
x42 vdd b3 net55 net48 b3b vss passtrans
x43 vdd b3b net53 net49 b3 vss passtrans
x44 vdd b3 net53 net50 b3b vss passtrans
x45 vdd b3b net54 net51 b3 vss passtrans
x46 vdd b3 net54 net52 b3b vss passtrans
x47 vdd vdd net61 net61 vss vss passtrans
.ends


* expanding   symbol:  passtrans.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rdac3v_8bit/xschem/passtrans.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rdac3v_8bit/xschem/passtrans.sch
.subckt passtrans vdd enab out in ena vss
*.PININFO enab:I ena:I vss:B vdd:B in:B out:B
XM1 in ena out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.65 nf=1 m=1
XM2 in enab out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends


* expanding   symbol:  rheo_level_shifter.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rheostat_8bit/xschem/rheo_level_shifter.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rheostat_8bit/xschem/rheo_level_shifter.sch
.subckt rheo_level_shifter avdd dvdd bit_out bitb_out bit_in dvss
*.PININFO bit_in:I bit_out:O bitb_out:O dvss:I dvdd:I avdd:I
x1 bit_in dvdd dvss dvss avdd avdd net1 sky130_fd_sc_hvl__lsbuflv2hv_1
x2 net1 dvss dvss avdd avdd net2 sky130_fd_sc_hvl__inv_2
x3 net2 dvss dvss avdd avdd net3 sky130_fd_sc_hvl__inv_4
x4 net3 dvss dvss avdd avdd bitb_out sky130_fd_sc_hvl__inv_8
x5 bitb_out dvss dvss avdd avdd bit_out sky130_fd_sc_hvl__inv_8
XXD1 dvss bit_in sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
.ends


* expanding   symbol:  rheo_column_dummy.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rheostat_8bit/xschem/rheo_column_dummy.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rheostat_8bit/xschem/rheo_column_dummy.sch
.subckt rheo_column_dummy vdd dum_in res_in res_out vss dum_out
*.PININFO res_in:B vss:B vdd:B dum_in:B res_out:B dum_out:B
x1 vdd vdd net17 net1 vss vss passtrans
x2 vdd vdd net16 net2 vss vss passtrans
x3 vdd vdd net15 net3 vss vss passtrans
x4 vdd vdd net14 net4 vss vss passtrans
x5 vdd vdd net13 net5 vss vss passtrans
x6 vdd vdd net12 net6 vss vss passtrans
x7 vdd vdd net10 net7 vss vss passtrans
x8 vdd vdd net11 res_in vss vss passtrans
x9 vdd vdd net8 dum_in vss vss passtrans
x10 vdd vdd net9 res_out vss vss passtrans
x11 vdd vdd net12 net12 vss vss passtrans
x12 vdd vdd net13 net13 vss vss passtrans
x13 vdd vdd net14 net14 vss vss passtrans
x14 vdd vdd net15 net15 vss vss passtrans
x15 vdd vdd net11 net11 vss vss passtrans
x16 vdd vdd net16 net16 vss vss passtrans
x17 vdd vdd net8 net8 vss vss passtrans
x18 vdd vdd net9 net9 vss vss passtrans
x19 vdd vdd net10 net10 vss vss passtrans
x20 vdd vdd net17 net17 vss vss passtrans
XR11 res_in dum_in sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR1 net7 res_in sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR2 net6 net7 sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR3 net5 net6 sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR4 net4 net5 sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR5 net3 net4 sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR6 net2 net3 sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR7 net1 net2 sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR8 res_out net1 sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR9 dum_out res_out sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
.ends


* expanding   symbol:  Stage0_clk_inv.sym # of pins=5
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_icrg_ip__ulpcomp/xschem/Stage0_clk_inv.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_icrg_ip__ulpcomp/xschem/Stage0_clk_inv.sch
.subckt Stage0_clk_inv dvddb clka clk clkb dvss
*.PININFO dvss:I dvddb:I clka:O clk:I clkb:O
XM22 clka clkb dvddb dvddb sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=1 m=1
XM8 clkb clk dvddb dvddb sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=1 m=1
XM6 clkb clk dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM21 clka clkb dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
.ends


* expanding   symbol:  Stage1.sym # of pins=10
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_icrg_ip__ulpcomp/xschem/Stage1.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_icrg_ip__ulpcomp/xschem/Stage1.sch
.subckt Stage1 avdd enab clka vinn vinp oneg opos avss dvss dvdd
*.PININFO avdd:I vinp:I vinn:I opos:O oneg:O clka:I enab:I dvdd:I avss:I dvss:I
XM1 net4 net5 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=2 m=2
x2 clka dvdd dvss dvss avdd avdd net2 sky130_fd_sc_hvl__lsbuflv2hv_1
XM6 net1 net2 net4 net4 sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=2 m=2
XM2 oneg vinp net1 net1 sky130_fd_pr__pfet_g5v0d10v5 L=1 W=20 nf=2 m=2
XM3 opos vinn net1 net1 sky130_fd_pr__pfet_g5v0d10v5 L=1 W=20 nf=2 m=2
XM4 net3 net3 avss avss sky130_fd_pr__nfet_03v3_nvt L=0.5 W=5 nf=1 m=2
XM8 opos net2 net3 net3 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM5 oneg net2 net3 net3 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
x1 enab dvdd dvss dvss avdd avdd net5 sky130_fd_sc_hvl__lsbuflv2hv_1
.ends


* expanding   symbol:  Stage2_latch.sym # of pins=8
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_icrg_ip__ulpcomp/xschem/Stage2_latch.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_icrg_ip__ulpcomp/xschem/Stage2_latch.sch
.subckt Stage2_latch dvdd enab dvddb clkb vout oneg opos dvss
*.PININFO clkb:I vout:O dvss:I dvdd:I opos:I oneg:I enab:I dvddb:O
XM18 vout net1 dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM19 vout net1 dvddb dvddb sky130_fd_pr__pfet_01v8 L=1 W=2 nf=1 m=1
XM15 net5 clkb dvss dvss sky130_fd_pr__nfet_03v3_nvt L=0.5 W=2 nf=1 m=1
XM9 net1 clkb dvddb dvddb sky130_fd_pr__pfet_01v8_hvt L=1 W=3 nf=1 m=2
XM10 net2 net1 dvddb dvddb sky130_fd_pr__pfet_01v8_hvt L=1 W=3 nf=1 m=2
XM11 net1 net2 dvddb dvddb sky130_fd_pr__pfet_01v8_hvt L=1 W=3 nf=1 m=2
XM12 net2 clkb dvddb dvddb sky130_fd_pr__pfet_01v8_hvt L=1 W=3 nf=1 m=2
XM1 dvddb enab dvdd dvdd sky130_fd_pr__pfet_01v8_hvt L=1 W=3 nf=1 m=2
XM2 net1 opos net3 dvss sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 m=1
XM3 net4 net1 net5 dvss sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 m=1
XM4 net3 net2 net5 dvss sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 m=1
XM5 net2 oneg net4 dvss sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 m=1
.ends


* expanding   symbol:  Stage0_ena_inv.sym # of pins=4
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_icrg_ip__ulpcomp/xschem/Stage0_ena_inv.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_icrg_ip__ulpcomp/xschem/Stage0_ena_inv.sch
.subckt Stage0_ena_inv dvdd ena enab dvss
*.PININFO ena:I dvdd:I dvss:I enab:O
XM25 enab ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=1 m=1
XM24 enab ena dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
.ends


* expanding   symbol:  buffer.sym # of pins=5
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_od_ip__tempsensor/xschem/buffer.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_od_ip__tempsensor/xschem/buffer.sch
.subckt buffer vdd vss vbias input output
*.PININFO output:O input:I vdd:I vss:I vbias:I
XM1 net2 input net1 vss sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
XM2 output output net1 vss sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
XM5 net1 vbias vss vss sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
XM4 output net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=10 W=1 nf=1 m=1
XM3 net2 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=10 W=1 nf=1 m=1
.ends


* expanding   symbol:  comp_hyst.sym # of pins=7
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_vbl_ip__overvoltage/xschem/comp_hyst.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_vbl_ip__overvoltage/xschem/comp_hyst.sch
.subckt comp_hyst dvdd out vref vin ena ibias dvss
*.PININFO dvdd:B vref:I vin:I out:O ibias:I ena:I dvss:B
XM5[0] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 m=1
XM5[1] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 m=1
XM3[0] net4 net4 dvdd dvdd sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 m=1
XM3[1] net4 net4 dvdd dvdd sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 m=1
XM7 net2 net4 dvdd dvdd sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 m=1
XM4[0] net3 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XM4[1] net3 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XM11 net5 net5 dvss dvss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 m=1
XM12 net1 net5 dvss dvss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 m=1
XM9 out net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=3 nf=1 m=1
XM10 out net2 dvss dvss sky130_fd_pr__nfet_01v8 L=1 W=3 nf=1 m=1
XM17 out ena_b dvss dvss sky130_fd_pr__nfet_01v8 L=3 W=1 nf=1 m=1
XM1[0] net4 vref net1 dvss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1.3 nf=1 m=1
XM1[1] net4 vref net1 dvss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1.3 nf=1 m=1
XM2[0] net3 vin net1 dvss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1.3 nf=1 m=1
XM2[1] net3 vin net1 dvss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1.3 nf=1 m=1
XM13 net5 ena_b dvss dvss sky130_fd_pr__nfet_01v8 L=3 W=1 nf=1 m=1
XM6[0] net4 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XM6[1] net4 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XM6[2] net4 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XM6[3] net4 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XM8 net2 net2 dvss dvss sky130_fd_pr__nfet_01v8 L=8 W=1 nf=1 m=1
XM16 net3 ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=3 W=1 nf=1 m=1
XM15 net4 ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=3 W=1 nf=1 m=1
XM14 net2 ena_b dvss dvss sky130_fd_pr__nfet_01v8 L=3 W=1 nf=1 m=1
XM18 ena_b ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=3 W=1 nf=1 m=1
XM19 ena_b ena dvss dvss sky130_fd_pr__nfet_01v8 L=3 W=1 nf=1 m=1
x1 ibias ena_b ena dvdd dvss net5 trans_gate
XMD16[0] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XMD16[1] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XMD16[2] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XMD16[3] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XMD16[4] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XMD16[5] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XMD8[0] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 m=1
XMD8[1] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 m=1
XMD1[0] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[1] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[2] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[3] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[4] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[5] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[6] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[7] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[8] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[9] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[10] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[11] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[12] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[13] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[14] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[15] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[16] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[17] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[18] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMD1[19] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XMDN8[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=1
XMDN8[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=1
XMDN1[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMDN1[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMDN1[2] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMDN1[3] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMDN2[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.3 nf=1 m=1
XMDN2[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.3 nf=1 m=1
XMDN2[2] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.3 nf=1 m=1
XMDN2[3] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.3 nf=1 m=1
XMDN2[4] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.3 nf=1 m=1
XMDN2[5] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.3 nf=1 m=1
XMDN2[6] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.3 nf=1 m=1
XMDN2[7] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1.3 nf=1 m=1
XD3 dvss vin sky130_fd_pr__diode_pw2nd_05v5 area=0.315e12 perim=2.3e6
XD1 dvss vref sky130_fd_pr__diode_pw2nd_05v5 area=0.315e12 perim=2.3e6
XD2 dvss ena sky130_fd_pr__diode_pw2nd_05v5 area=0.315e12 perim=2.3e6
.ends


* expanding   symbol:  ov_multiplexer.sym # of pins=27
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_vbl_ip__overvoltage/xschem/ov_multiplexer.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_vbl_ip__overvoltage/xschem/ov_multiplexer.sch
.subckt ov_multiplexer in_0000 in_0001 in_0010 in_0011 in_0100 in_0101 in_0110 avdd vss in_0111 vtrip_3 vtrip_3_b vtrip_2
+ vtrip_2_b vtrip_1 out vtrip_1_b vtrip_0 vtrip_0_b in_1000 in_1001 in_1010 in_1011 in_1100 in_1101 in_1110 in_1111
*.PININFO in_0000:I in_0001:I in_0010:I in_0011:I in_0100:I in_0101:I in_0110:I in_0111:I in_1000:I in_1001:I in_1010:I in_1011:I
*+ in_1110:I in_1111:I in_1100:I in_1101:I out:O vtrip_3:I vtrip_3_b:I vtrip_2:I vtrip_2_b:I vtrip_1:I vtrip_1_b:I vtrip_0:I vtrip_0_b:I
*+ avdd:B vss:B
x1 net5 vtrip_3 vtrip_3_b avdd vss out trans_gate_mux
x2 net6 vtrip_3_b vtrip_3 avdd vss out trans_gate_mux
x3 net2 vtrip_2 vtrip_2_b avdd vss net6 trans_gate_mux
x4 net4 vtrip_2_b vtrip_2 avdd vss net5 trans_gate_mux
x5 net3 vtrip_2_b vtrip_2 avdd vss net6 trans_gate_mux
x6 net1 vtrip_2 vtrip_2_b avdd vss net5 trans_gate_mux
x7 net7 vtrip_1 vtrip_1_b avdd vss net1 trans_gate_mux
x8 net8 vtrip_1_b vtrip_1 avdd vss net1 trans_gate_mux
x9 net9 vtrip_1 vtrip_1_b avdd vss net4 trans_gate_mux
x10 net10 vtrip_1_b vtrip_1 avdd vss net4 trans_gate_mux
x11 net11 vtrip_1 vtrip_1_b avdd vss net2 trans_gate_mux
x12 net12 vtrip_1_b vtrip_1 avdd vss net2 trans_gate_mux
x13 net13 vtrip_1 vtrip_1_b avdd vss net3 trans_gate_mux
x14 net14 vtrip_1_b vtrip_1 avdd vss net3 trans_gate_mux
x15 in_0000 vtrip_0 vtrip_0_b avdd vss net7 trans_gate_mux
x16 in_0001 vtrip_0_b vtrip_0 avdd vss net7 trans_gate_mux
x17 in_0010 vtrip_0 vtrip_0_b avdd vss net8 trans_gate_mux
x18 in_0011 vtrip_0_b vtrip_0 avdd vss net8 trans_gate_mux
x19 in_0100 vtrip_0 vtrip_0_b avdd vss net9 trans_gate_mux
x20 in_0101 vtrip_0_b vtrip_0 avdd vss net9 trans_gate_mux
x21 in_0110 vtrip_0 vtrip_0_b avdd vss net10 trans_gate_mux
x22 in_0111 vtrip_0_b vtrip_0 avdd vss net10 trans_gate_mux
x23 in_1000 vtrip_0 vtrip_0_b avdd vss net11 trans_gate_mux
x24 in_1001 vtrip_0_b vtrip_0 avdd vss net11 trans_gate_mux
x25 in_1010 vtrip_0 vtrip_0_b avdd vss net12 trans_gate_mux
x26 in_1011 vtrip_0_b vtrip_0 avdd vss net12 trans_gate_mux
x27 in_1100 vtrip_0 vtrip_0_b avdd vss net13 trans_gate_mux
x28 in_1101 vtrip_0_b vtrip_0 avdd vss net13 trans_gate_mux
x29 in_1110 vtrip_0 vtrip_0_b avdd vss net14 trans_gate_mux
x30 in_1111 vtrip_0_b vtrip_0 avdd vss net14 trans_gate_mux
XD1 vss vtrip_0 sky130_fd_pr__diode_pw2nd_05v5 area=3.15e11 perim=2.3e6
XD2 vss vtrip_0 sky130_fd_pr__diode_pw2nd_05v5 area=3.15e11 perim=2.3e6
XD3 vss vtrip_0_b sky130_fd_pr__diode_pw2nd_05v5 area=3.15e11 perim=2.3e6
XD4 vss vtrip_0_b sky130_fd_pr__diode_pw2nd_05v5 area=3.15e11 perim=2.3e6
XD5 vss vtrip_1 sky130_fd_pr__diode_pw2nd_05v5 area=3.15e11 perim=2.3e6
XD6 vss vtrip_1 sky130_fd_pr__diode_pw2nd_05v5 area=3.15e11 perim=2.3e6
XD7 vss vtrip_1_b sky130_fd_pr__diode_pw2nd_05v5 area=3.15e11 perim=2.3e6
XD8 vss vtrip_1_b sky130_fd_pr__diode_pw2nd_05v5 area=3.15e11 perim=2.3e6
XD9 vss vtrip_2 sky130_fd_pr__diode_pw2nd_05v5 area=3.15e11 perim=2.3e6
XD11 vss vtrip_2_b sky130_fd_pr__diode_pw2nd_05v5 area=3.15e11 perim=2.3e6
XD10 vss vtrip_3 sky130_fd_pr__diode_pw2nd_05v5 area=3.15e11 perim=2.3e6
XD12 vss vtrip_3_b sky130_fd_pr__diode_pw2nd_05v5 area=3.15e11 perim=2.3e6
.ends


* expanding   symbol:  ov_voltage_divider.sym # of pins=19
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_vbl_ip__overvoltage/xschem/ov_voltage_divider.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_vbl_ip__overvoltage/xschem/ov_voltage_divider.sch
.subckt ov_voltage_divider avdd out_0000 out_0001 out_0010 out_0011 out_0100 out_0101 out_0110 out_0111 out_1000 out_1001 out_1010
+ out_1011 out_1100 out_1101 out_1110 out_1111 avss ena
*.PININFO ena:I avss:B avdd:B out_1111:O out_1110:O out_1101:O out_1100:O out_1011:O out_1010:O out_1001:O out_1000:O out_0111:O
*+ out_0110:O out_0101:O out_0100:O out_0011:O out_0010:O out_0001:O out_0000:O
XM1 res[0] ena avss avss sky130_fd_pr__nfet_g5v0d10v5 L=3 W=3 nf=1 m=1
XRA[28] res[28] res[29] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[27] res[27] res[28] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[26] res[26] res[27] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[25] res[25] res[26] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[24] res[24] res[25] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[23] res[23] res[24] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[22] res[22] res[23] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[21] res[21] res[22] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[20] res[20] res[21] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[19] res[19] res[20] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[18] res[18] res[19] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[17] res[17] res[18] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[16] res[16] res[17] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[15] res[15] res[16] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[14] res[14] res[15] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[13] res[13] res[14] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[12] res[12] res[13] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[11] res[11] res[12] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[10] res[10] res[11] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[9] res[9] res[10] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[8] res[8] res[9] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[7] res[7] res[8] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[6] res[6] res[7] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[5] res[5] res[6] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[4] res[4] res[5] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[3] res[3] res[4] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[2] res[2] res[3] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[1] res[1] res[2] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRA[0] res[0] res[1] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR1 res[29] out_1111 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR2 out_1111 out_1110 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR3 out_1110 out_1101 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR4 out_1101 out_1100 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR5 out_1100 out_1011 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR6 out_1011 out_1010 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR7 out_1010 out_1001 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR8 out_1001 out_1000 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR9 out_1000 out_0111 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR10 out_0111 net1 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR11 net1 out_0110 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR12 out_0110 out_0101 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR13 out_0101 net2 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR14 net2 out_0100 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR15 out_0100 out_0011 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR16 out_0011 net3 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR17 net3 out_0010 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR18 out_0010 net4 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR19 net4 out_0001 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR20 out_0001 net5 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR21 net5 out_0000 avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR22 out_0000 res[30] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[85] res[115] res[116] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[84] res[114] res[115] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[83] res[113] res[114] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[82] res[112] res[113] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[81] res[111] res[112] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[80] res[110] res[111] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[79] res[109] res[110] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[78] res[108] res[109] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[77] res[107] res[108] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[76] res[106] res[107] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[75] res[105] res[106] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[74] res[104] res[105] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[73] res[103] res[104] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[72] res[102] res[103] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[71] res[101] res[102] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[70] res[100] res[101] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[69] res[99] res[100] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[68] res[98] res[99] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[67] res[97] res[98] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[66] res[96] res[97] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[65] res[95] res[96] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[64] res[94] res[95] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[63] res[93] res[94] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[62] res[92] res[93] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[61] res[91] res[92] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[60] res[90] res[91] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[59] res[89] res[90] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[58] res[88] res[89] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[57] res[87] res[88] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[56] res[86] res[87] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[55] res[85] res[86] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[54] res[84] res[85] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[53] res[83] res[84] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[52] res[82] res[83] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[51] res[81] res[82] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[50] res[80] res[81] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[49] res[79] res[80] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[48] res[78] res[79] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[47] res[77] res[78] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[46] res[76] res[77] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[45] res[75] res[76] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[44] res[74] res[75] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[43] res[73] res[74] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[42] res[72] res[73] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[41] res[71] res[72] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[40] res[70] res[71] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[39] res[69] res[70] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[38] res[68] res[69] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[37] res[67] res[68] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[36] res[66] res[67] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[35] res[65] res[66] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[34] res[64] res[65] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[33] res[63] res[64] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[32] res[62] res[63] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[31] res[61] res[62] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[30] res[60] res[61] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[29] res[59] res[60] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[28] res[58] res[59] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[27] res[57] res[58] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[26] res[56] res[57] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[25] res[55] res[56] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[24] res[54] res[55] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[23] res[53] res[54] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[22] res[52] res[53] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[21] res[51] res[52] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[20] res[50] res[51] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[19] res[49] res[50] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[18] res[48] res[49] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[17] res[47] res[48] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[16] res[46] res[47] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[15] res[45] res[46] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[14] res[44] res[45] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[13] res[43] res[44] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[12] res[42] res[43] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[11] res[41] res[42] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[10] res[40] res[41] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[9] res[39] res[40] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[8] res[38] res[39] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[7] res[37] res[38] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[6] res[36] res[37] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[5] res[35] res[36] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[4] res[34] res[35] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[3] res[33] res[34] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[2] res[32] res[33] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[1] res[31] res[32] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRB[0] res[30] res[31] avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XR23 res[116] avdd avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=1 m=1
XRdummy1 avss avss avss sky130_fd_pr__res_xhigh_po_1p41 L=14.1 mult=6 m=6
XRdummy2 avss avss avss sky130_fd_pr__res_xhigh_po_1p41 L=1.41 mult=96 m=96
XD1 avss ena sky130_fd_pr__diode_pw2nd_05v5 area=3.15e11 perim=2.3e6
.ends


* expanding   symbol:  ov_level_shifter.sym # of pins=7
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_vbl_ip__overvoltage/xschem/ov_level_shifter.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_vbl_ip__overvoltage/xschem/ov_level_shifter.sch
.subckt ov_level_shifter avdd dvdd in out out_b avss dvss
*.PININFO avdd:B out_b:O out:O avss:B dvdd:B in:I dvss:B
XM1 in_b in dvss dvss sky130_fd_pr__nfet_01v8 L=3 W=1 nf=1 m=1
XM2 in_b in dvdd dvdd sky130_fd_pr__pfet_01v8 L=3 W=1 nf=1 m=1
XM3 out_b out avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1 nf=1 m=1
XM4 out out_b avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1 nf=1 m=1
XM8 out in_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=3 W=2 nf=1 m=1
XM7 out_b in avss avss sky130_fd_pr__nfet_g5v0d10v5 L=3 W=2 nf=1 m=1
XD3 dvss in sky130_fd_pr__diode_pw2nd_05v5 area=0.315e12 perim=2.3e6
.ends


* expanding   symbol:  dac_half.sym # of pins=21
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rdac3v_8bit/xschem/dac_half.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rdac3v_8bit/xschem/dac_half.sch
.subckt dac_half vdd vss b3 b4 b3b b4b b5 res_in b6 b0 dum_in b6b b5b b0b b1 b1b b2 b2b out res_out dum_out
*.PININFO res_in:B res_out:B out:B vdd:B vss:B b3:I b3b:I b5:I b5b:I b6:I b6b:I dum_out:B dum_in:B b4:I b4b:I b0:I b0b:I b1:I
*+ b1b:I b2:I b2b:I
x1 b2 b2b b1 b1b b0 b0b vdd net9 net8 net44 net16 vss net15 dac_column
x2 b2 b2b b1 b1b b0 b0b vdd net10 net7 net43 net8 vss net9 dac_column
x3 b2 b2b b1 b1b b0 b0b vdd net11 net6 net42 net7 vss net10 dac_column
x4 b2 b2b b1 b1b b0 b0b vdd net12 net5 net41 net6 vss net11 dac_column
x5 b2 b2b b1 b1b b0 b0b vdd net13 net4 net40 net5 vss net12 dac_column
x6 b2 b2b b1 b1b b0 b0b vdd net14 net3 net39 net4 vss net13 dac_column
x7 b2 b2b b1 b1b b0 b0b vdd net2 net1 net38 net3 vss net14 dac_column
x8 b2 b2b b1 b1b b0 b0b vdd dum_in res_in net37 net1 vss net2 dac_column
x9 b2 b2b b1 b1b b0 b0b vdd net25 net24 net52 res_out vss dum_out dac_column
x10 b2 b2b b1 b1b b0 b0b vdd net26 net23 net51 net24 vss net25 dac_column
x11 b2 b2b b1 b1b b0 b0b vdd net27 net22 net50 net23 vss net26 dac_column
x12 b2 b2b b1 b1b b0 b0b vdd net28 net21 net49 net22 vss net27 dac_column
x13 b2 b2b b1 b1b b0 b0b vdd net29 net20 net48 net21 vss net28 dac_column
x14 b2 b2b b1 b1b b0 b0b vdd net30 net19 net47 net20 vss net29 dac_column
x15 b2 b2b b1 b1b b0 b0b vdd net18 net17 net46 net19 vss net30 dac_column
x16 b2 b2b b1 b1b b0 b0b vdd net15 net16 net45 net17 vss net18 dac_column
x17 vdd b4 net31 net54 b4b vss passtrans
x18 vdd b4b net31 net53 b4 vss passtrans
x19 vdd b4 net32 net55 b4b vss passtrans
x20 vdd b4b net32 net56 b4 vss passtrans
x21 vdd b4 net33 net57 b4b vss passtrans
x22 vdd b4b net33 net58 b4 vss passtrans
x23 vdd b4 net34 net59 b4b vss passtrans
x24 vdd b4b net34 net60 b4 vss passtrans
x25 vdd b5b net36 net34 b5 vss passtrans
x26 vdd b5 net36 net33 b5b vss passtrans
x27 vdd b5b net35 net32 b5 vss passtrans
x28 vdd b5 net35 net31 b5b vss passtrans
x29 vdd b6b out net36 b6 vss passtrans
x30 vdd b6 out net35 b6b vss passtrans
x33 vdd b3b net60 net37 b3 vss passtrans
x31 vdd b3 net60 net38 b3b vss passtrans
x32 vdd b3b net59 net39 b3 vss passtrans
x34 vdd b3 net59 net40 b3b vss passtrans
x35 vdd b3b net58 net41 b3 vss passtrans
x36 vdd b3 net58 net42 b3b vss passtrans
x37 vdd b3b net57 net43 b3 vss passtrans
x38 vdd b3 net57 net44 b3b vss passtrans
x39 vdd b3b net56 net45 b3 vss passtrans
x40 vdd b3 net56 net46 b3b vss passtrans
x41 vdd b3b net55 net47 b3 vss passtrans
x42 vdd b3 net55 net48 b3b vss passtrans
x43 vdd b3b net53 net49 b3 vss passtrans
x44 vdd b3 net53 net50 b3b vss passtrans
x45 vdd b3b net54 net51 b3 vss passtrans
x46 vdd b3 net54 net52 b3b vss passtrans
x47 vdd vdd net61 net61 vss vss passtrans
.ends


* expanding   symbol:  level_shifter.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rdac3v_8bit/xschem/level_shifter.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rdac3v_8bit/xschem/level_shifter.sch
.subckt level_shifter vdd dvdd bit_out bitb_out bit_in dvss
*.PININFO bit_in:I bit_out:O bitb_out:O dvss:I dvdd:I vdd:I
x1 bit_in dvdd dvss dvss vdd vdd net1 sky130_fd_sc_hvl__lsbuflv2hv_1
x2 net1 dvss dvss vdd vdd net2 sky130_fd_sc_hvl__inv_2
x3 net2 dvss dvss vdd vdd net3 sky130_fd_sc_hvl__inv_4
x4 net3 dvss dvss vdd vdd bitb_out sky130_fd_sc_hvl__inv_8
x5 bitb_out dvss dvss vdd vdd bit_out sky130_fd_sc_hvl__inv_8
XXD1 dvss bit_in sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
.ends


* expanding   symbol:  dac_column_dummy.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rdac3v_8bit/xschem/dac_column_dummy.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rdac3v_8bit/xschem/dac_column_dummy.sch
.subckt dac_column_dummy vdd dum_in res_in res_out vss dum_out
*.PININFO res_in:B vss:B vdd:B dum_in:B res_out:B dum_out:B
x1 vdd vdd net17 net1 vss vss passtrans
XR1 res_out net1 vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
x2 vdd vdd net16 net2 vss vss passtrans
x3 vdd vdd net15 net3 vss vss passtrans
x4 vdd vdd net14 net4 vss vss passtrans
x5 vdd vdd net13 net5 vss vss passtrans
x6 vdd vdd net12 net6 vss vss passtrans
x7 vdd vdd net10 net7 vss vss passtrans
x8 vdd vdd net11 res_in vss vss passtrans
x9 vdd vdd net8 dum_in vss vss passtrans
x10 vdd vdd net9 res_out vss vss passtrans
XR2 net1 net2 vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR3 net2 net3 vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR4 net3 net4 vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR5 net4 net5 vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR6 net5 net6 vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR7 net6 net7 vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR9 net7 res_in vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR10 res_in dum_in vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR12 dum_out res_out vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
x11 vdd vdd net12 net12 vss vss passtrans
x12 vdd vdd net13 net13 vss vss passtrans
x13 vdd vdd net14 net14 vss vss passtrans
x14 vdd vdd net15 net15 vss vss passtrans
x15 vdd vdd net11 net11 vss vss passtrans
x16 vdd vdd net16 net16 vss vss passtrans
x17 vdd vdd net8 net8 vss vss passtrans
x18 vdd vdd net9 net9 vss vss passtrans
x19 vdd vdd net10 net10 vss vss passtrans
x20 vdd vdd net17 net17 vss vss passtrans
.ends


* expanding   symbol:  follower_amp.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rdac3v_8bit/dependencies/sky130_ef_ip__samplehold/xschem/follower_amp.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rdac3v_8bit/dependencies/sky130_ef_ip__samplehold/xschem/follower_amp.sch
.subckt follower_amp vdd out ena vss in vsub
*.PININFO in:I vdd:I vss:I out:O ena:I vsub:I
XM4 pdrv1 net1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM5 vdd net1 net1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM10 vss nbias nbias vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=4 m=1
XM20 out pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=280 nf=280 m=1
XM22 out ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=4 m=1
XM24 pbias nbias vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM25 vdd pbias pbias vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM26 vcomp pbias vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM27 net2 out vcomp vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM28 vcomp in ndrv vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM29 ndrv net2 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM30 vss net2 net2 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM1 net1 out vcomn1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM2 vcomn1 in pdrv1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM3 pdrv2 net3 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM6 vdd net3 net3 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM7 vcomn2 nbias vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM12 vdd pdrv2 out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=20 nf=20 m=1
XXD1 vss in sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
XM13 net4 ena nbias vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XXD2 vss ena sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
XM11 pdrv2 in vcomn2 vss sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 m=1
XM9 net3 out vcomn2 vss sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 m=1
XM8 vcomn1 nbias vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XR2 net4 vdd vss sky130_fd_pr__res_xhigh_po_0p35 L=35 mult=1 m=1
.ends


* expanding   symbol:  isolated_switch_large.sym # of pins=8
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/isolated_switch_large.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/isolated_switch_large.sch
.subckt isolated_switch_large avss on out in avdd dvdd dvss off
*.PININFO on:I avss:B out:B in:B avdd:B dvdd:B dvss:B off:I
x2 on dvdd dvss dvss avdd avdd net1 sky130_fd_sc_hvl__lsbuflv2hv_1
x1 net1 net2 avss out in avdd net3 isolated_switch_3
x3 off dvdd dvss dvss avdd avdd net3 sky130_fd_sc_hvl__lsbuflv2hv_1
x4 net1 dvss dvss avdd avdd net2 sky130_fd_sc_hvl__inv_1
x5 on dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x6 off dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
.ends


* expanding   symbol:  isolated_switch_xlarge.sym # of pins=8
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/isolated_switch_xlarge.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/isolated_switch_xlarge.sch
.subckt isolated_switch_xlarge avss on out in avdd dvdd dvss off
*.PININFO on:I avss:B out:B in:B avdd:B dvdd:B dvss:B off:I
x2 on dvdd dvss dvss avdd avdd net1 sky130_fd_sc_hvl__lsbuflv2hv_1
x1 net1 net2 avss out in avdd net3 isolated_switch_4
x3 off dvdd dvss dvss avdd avdd net3 sky130_fd_sc_hvl__lsbuflv2hv_1
x4 net1 dvss dvss avdd avdd net2 sky130_fd_sc_hvl__inv_1
x5 on dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x6 off dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
.ends


* expanding   symbol:  simplest_analog_switch_ena1v8.sym # of pins=7
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/simplest_analog_switch_ena1v8.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/simplest_analog_switch_ena1v8.sch
.subckt simplest_analog_switch_ena1v8 avss on out in avdd dvdd dvss
*.PININFO on:I avss:B out:B in:B avdd:B dvdd:B dvss:B
x2 on dvdd dvss dvss avdd avdd net3 sky130_fd_sc_hvl__lsbuflv2hv_1
x3 net1 net2 avss out in avdd simple_analog_switch_2
x1 net3 dvss dvss avdd avdd net2 sky130_fd_sc_hvl__inv_2
x4 net2 dvss dvss avdd avdd net1 sky130_fd_sc_hvl__inv_2
x5[1] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x5[0] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x5 on dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
.ends


* expanding   symbol:  simple_analog_switch_2.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch_2.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch_2.sch
.subckt simple_analog_switch_2 on off vss out in vdd
*.PININFO on:I out:B vdd:B vss:B in:B off:I
XM1 in on out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 nf=4 m=1
XM2 in off out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=40 nf=8 m=1
.ends


* expanding   symbol:  bias_generator_fe.sym # of pins=15
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/bias_generator_fe.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/bias_generator_fe.sch
.subckt bias_generator_fe avdd ena vbg src_test0 avss dvdd ena_src_test0 ref_sel_vbg ref_in dvss nbias pcasc pbias snk_test0
+ ena_snk_test0
*.PININFO ref_in:I avss:B ref_sel_vbg:I avdd:B ena_src_test0:I ena_snk_test0:I src_test0:B snk_test0:B vbg:I ena:I dvdd:B dvss:B
*+ pcasc:O pbias:O nbias:O
x2[19] net1 ena_3v3 nbias nbias avss bias_nstack
x2[18] net1 ena_3v3 nbias nbias avss bias_nstack
x2[17] net1 ena_3v3 nbias nbias avss bias_nstack
x2[16] net1 ena_3v3 nbias nbias avss bias_nstack
x2[15] net1 ena_3v3 nbias nbias avss bias_nstack
x2[14] net1 ena_3v3 nbias nbias avss bias_nstack
x2[13] net1 ena_3v3 nbias nbias avss bias_nstack
x2[12] net1 ena_3v3 nbias nbias avss bias_nstack
x2[11] net1 ena_3v3 nbias nbias avss bias_nstack
x2[10] net1 ena_3v3 nbias nbias avss bias_nstack
x2[9] net1 ena_3v3 nbias nbias avss bias_nstack
x2[8] net1 ena_3v3 nbias nbias avss bias_nstack
x2[7] net1 ena_3v3 nbias nbias avss bias_nstack
x2[6] net1 ena_3v3 nbias nbias avss bias_nstack
x2[5] net1 ena_3v3 nbias nbias avss bias_nstack
x2[4] net1 ena_3v3 nbias nbias avss bias_nstack
x2[3] net1 ena_3v3 nbias nbias avss bias_nstack
x2[2] net1 ena_3v3 nbias nbias avss bias_nstack
x2[1] net1 ena_3v3 nbias nbias avss bias_nstack
x2[0] net1 ena_3v3 nbias nbias avss bias_nstack
XR4 pcasc ref_in avss sky130_fd_pr__res_high_po_0p35 L=1500 mult=1 m=1
x4 pbias enb_vbg_3v3 net2 nbias avss bias_nstack
x2 avdd pbias pcasc net5 ena_vbg_3v3 avss pbias bias_pstack
x13[9] avdd pbias pcasc net6[9] enb_test0_3v3 avss src_test0 bias_pstack
x13[8] avdd pbias pcasc net6[8] enb_test0_3v3 avss src_test0 bias_pstack
x13[7] avdd pbias pcasc net6[7] enb_test0_3v3 avss src_test0 bias_pstack
x13[6] avdd pbias pcasc net6[6] enb_test0_3v3 avss src_test0 bias_pstack
x13[5] avdd pbias pcasc net6[5] enb_test0_3v3 avss src_test0 bias_pstack
x13[4] avdd pbias pcasc net6[4] enb_test0_3v3 avss src_test0 bias_pstack
x13[3] avdd pbias pcasc net6[3] enb_test0_3v3 avss src_test0 bias_pstack
x13[2] avdd pbias pcasc net6[2] enb_test0_3v3 avss src_test0 bias_pstack
x13[1] avdd pbias pcasc net6[1] enb_test0_3v3 avss src_test0 bias_pstack
x13[0] avdd pbias pcasc net6[0] enb_test0_3v3 avss src_test0 bias_pstack
x17[1] snk_test0 ena_test0_3v3 net7[1] nbias avss bias_nstack
x17[0] snk_test0 ena_test0_3v3 net7[0] nbias avss bias_nstack
x1 ref_sel_vbg dvdd dvss dvss avdd avdd ena_vbg_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x11 ena_snk_test0 dvdd dvss dvss avdd avdd ena_test0_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x23 ena_src_test0 dvdd dvss dvss avdd avdd net4 sky130_fd_sc_hvl__lsbuflv2hv_1
x24 ena_vbg_3v3 dvss dvss avdd avdd enb_vbg_3v3 sky130_fd_sc_hvl__inv_2
x35 net4 dvss dvss avdd avdd enb_test0_3v3 sky130_fd_sc_hvl__inv_2
x3 avdd pbias vbg vfb nbias avss ena_vbg_3v3 bias_amp
XR1 avss net3 avss sky130_fd_pr__res_high_po_0p35 L=2008 mult=1 m=1
XC1 pbias vfb sky130_fd_pr__cap_mim_m3_1 W=5 L=5 m=8
x36 ena dvdd dvss dvss avdd avdd ena_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
* noconn #net2
* noconn #net7
* noconn #net6
XR2 net1 pcasc avss sky130_fd_pr__res_high_po_0p35 L=900 mult=1 m=1
Vmeas vfb net3 0
.save i(vmeas)
x19[11] avdd pbias pcasc net8[11] enb_vbg_3v3 avss vfb bias_pstack
x19[10] avdd pbias pcasc net8[10] enb_vbg_3v3 avss vfb bias_pstack
x19[9] avdd pbias pcasc net8[9] enb_vbg_3v3 avss vfb bias_pstack
x19[8] avdd pbias pcasc net8[8] enb_vbg_3v3 avss vfb bias_pstack
x19[7] avdd pbias pcasc net8[7] enb_vbg_3v3 avss vfb bias_pstack
x19[6] avdd pbias pcasc net8[6] enb_vbg_3v3 avss vfb bias_pstack
x19[5] avdd pbias pcasc net8[5] enb_vbg_3v3 avss vfb bias_pstack
x19[4] avdd pbias pcasc net8[4] enb_vbg_3v3 avss vfb bias_pstack
x19[3] avdd pbias pcasc net8[3] enb_vbg_3v3 avss vfb bias_pstack
x19[2] avdd pbias pcasc net8[2] enb_vbg_3v3 avss vfb bias_pstack
x19[1] avdd pbias pcasc net8[1] enb_vbg_3v3 avss vfb bias_pstack
x19[0] avdd pbias pcasc net8[0] enb_vbg_3v3 avss vfb bias_pstack
* noconn #net8
* noconn #net5
XD1 avss vbg sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
x5[1] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x5[0] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x5 ref_sel_vbg dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x6 ena dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x7 ena_src_test0 dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x8 ena_snk_test0 dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
.ends


* expanding   symbol:  bias_generator_idac_be.sym # of pins=10
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/bias_generator_idac_be.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/bias_generator_idac_be.sch
.subckt bias_generator_idac_be dvdd dvss ena[7] ena[6] ena[5] ena[4] ena[3] ena[2] ena[1] ena[0] avdd pcasc pbias src_out snk_out
+ nbias avss
*.PININFO avss:B avdd:B src_out:B ena[7:0]:I dvdd:B dvss:B pcasc:I pbias:I nbias:I snk_out:B
x3 snk_out avss net1 nbias avss bias_nstack
x1 avdd pbias pcasc net2 avdd avss src_out bias_pstack
x8 avdd pbias pcasc net3 enb_bit0 avss src_out bias_pstack
x4[1] avdd pbias pcasc net4[1] enb_bit1 avss src_out bias_pstack
x4[0] avdd pbias pcasc net4[0] enb_bit1 avss src_out bias_pstack
x5[3] avdd pbias pcasc net5[3] enb_bit2 avss src_out bias_pstack
x5[2] avdd pbias pcasc net5[2] enb_bit2 avss src_out bias_pstack
x5[1] avdd pbias pcasc net5[1] enb_bit2 avss src_out bias_pstack
x5[0] avdd pbias pcasc net5[0] enb_bit2 avss src_out bias_pstack
x6[7] avdd pbias pcasc net6[7] enb_bit3 avss src_out bias_pstack
x6[6] avdd pbias pcasc net6[6] enb_bit3 avss src_out bias_pstack
x6[5] avdd pbias pcasc net6[5] enb_bit3 avss src_out bias_pstack
x6[4] avdd pbias pcasc net6[4] enb_bit3 avss src_out bias_pstack
x6[3] avdd pbias pcasc net6[3] enb_bit3 avss src_out bias_pstack
x6[2] avdd pbias pcasc net6[2] enb_bit3 avss src_out bias_pstack
x6[1] avdd pbias pcasc net6[1] enb_bit3 avss src_out bias_pstack
x6[0] avdd pbias pcasc net6[0] enb_bit3 avss src_out bias_pstack
x7[15] avdd pbias pcasc net7[15] enb_bit4 avss src_out bias_pstack
x7[14] avdd pbias pcasc net7[14] enb_bit4 avss src_out bias_pstack
x7[13] avdd pbias pcasc net7[13] enb_bit4 avss src_out bias_pstack
x7[12] avdd pbias pcasc net7[12] enb_bit4 avss src_out bias_pstack
x7[11] avdd pbias pcasc net7[11] enb_bit4 avss src_out bias_pstack
x7[10] avdd pbias pcasc net7[10] enb_bit4 avss src_out bias_pstack
x7[9] avdd pbias pcasc net7[9] enb_bit4 avss src_out bias_pstack
x7[8] avdd pbias pcasc net7[8] enb_bit4 avss src_out bias_pstack
x7[7] avdd pbias pcasc net7[7] enb_bit4 avss src_out bias_pstack
x7[6] avdd pbias pcasc net7[6] enb_bit4 avss src_out bias_pstack
x7[5] avdd pbias pcasc net7[5] enb_bit4 avss src_out bias_pstack
x7[4] avdd pbias pcasc net7[4] enb_bit4 avss src_out bias_pstack
x7[3] avdd pbias pcasc net7[3] enb_bit4 avss src_out bias_pstack
x7[2] avdd pbias pcasc net7[2] enb_bit4 avss src_out bias_pstack
x7[1] avdd pbias pcasc net7[1] enb_bit4 avss src_out bias_pstack
x7[0] avdd pbias pcasc net7[0] enb_bit4 avss src_out bias_pstack
x11[31] avdd pbias pcasc net8[31] enb_bit5 avss src_out bias_pstack
x11[30] avdd pbias pcasc net8[30] enb_bit5 avss src_out bias_pstack
x11[29] avdd pbias pcasc net8[29] enb_bit5 avss src_out bias_pstack
x11[28] avdd pbias pcasc net8[28] enb_bit5 avss src_out bias_pstack
x11[27] avdd pbias pcasc net8[27] enb_bit5 avss src_out bias_pstack
x11[26] avdd pbias pcasc net8[26] enb_bit5 avss src_out bias_pstack
x11[25] avdd pbias pcasc net8[25] enb_bit5 avss src_out bias_pstack
x11[24] avdd pbias pcasc net8[24] enb_bit5 avss src_out bias_pstack
x11[23] avdd pbias pcasc net8[23] enb_bit5 avss src_out bias_pstack
x11[22] avdd pbias pcasc net8[22] enb_bit5 avss src_out bias_pstack
x11[21] avdd pbias pcasc net8[21] enb_bit5 avss src_out bias_pstack
x11[20] avdd pbias pcasc net8[20] enb_bit5 avss src_out bias_pstack
x11[19] avdd pbias pcasc net8[19] enb_bit5 avss src_out bias_pstack
x11[18] avdd pbias pcasc net8[18] enb_bit5 avss src_out bias_pstack
x11[17] avdd pbias pcasc net8[17] enb_bit5 avss src_out bias_pstack
x11[16] avdd pbias pcasc net8[16] enb_bit5 avss src_out bias_pstack
x11[15] avdd pbias pcasc net8[15] enb_bit5 avss src_out bias_pstack
x11[14] avdd pbias pcasc net8[14] enb_bit5 avss src_out bias_pstack
x11[13] avdd pbias pcasc net8[13] enb_bit5 avss src_out bias_pstack
x11[12] avdd pbias pcasc net8[12] enb_bit5 avss src_out bias_pstack
x11[11] avdd pbias pcasc net8[11] enb_bit5 avss src_out bias_pstack
x11[10] avdd pbias pcasc net8[10] enb_bit5 avss src_out bias_pstack
x11[9] avdd pbias pcasc net8[9] enb_bit5 avss src_out bias_pstack
x11[8] avdd pbias pcasc net8[8] enb_bit5 avss src_out bias_pstack
x11[7] avdd pbias pcasc net8[7] enb_bit5 avss src_out bias_pstack
x11[6] avdd pbias pcasc net8[6] enb_bit5 avss src_out bias_pstack
x11[5] avdd pbias pcasc net8[5] enb_bit5 avss src_out bias_pstack
x11[4] avdd pbias pcasc net8[4] enb_bit5 avss src_out bias_pstack
x11[3] avdd pbias pcasc net8[3] enb_bit5 avss src_out bias_pstack
x11[2] avdd pbias pcasc net8[2] enb_bit5 avss src_out bias_pstack
x11[1] avdd pbias pcasc net8[1] enb_bit5 avss src_out bias_pstack
x11[0] avdd pbias pcasc net8[0] enb_bit5 avss src_out bias_pstack
x12[63] avdd pbias pcasc net9[63] enb_bit6 avss src_out bias_pstack
x12[62] avdd pbias pcasc net9[62] enb_bit6 avss src_out bias_pstack
x12[61] avdd pbias pcasc net9[61] enb_bit6 avss src_out bias_pstack
x12[60] avdd pbias pcasc net9[60] enb_bit6 avss src_out bias_pstack
x12[59] avdd pbias pcasc net9[59] enb_bit6 avss src_out bias_pstack
x12[58] avdd pbias pcasc net9[58] enb_bit6 avss src_out bias_pstack
x12[57] avdd pbias pcasc net9[57] enb_bit6 avss src_out bias_pstack
x12[56] avdd pbias pcasc net9[56] enb_bit6 avss src_out bias_pstack
x12[55] avdd pbias pcasc net9[55] enb_bit6 avss src_out bias_pstack
x12[54] avdd pbias pcasc net9[54] enb_bit6 avss src_out bias_pstack
x12[53] avdd pbias pcasc net9[53] enb_bit6 avss src_out bias_pstack
x12[52] avdd pbias pcasc net9[52] enb_bit6 avss src_out bias_pstack
x12[51] avdd pbias pcasc net9[51] enb_bit6 avss src_out bias_pstack
x12[50] avdd pbias pcasc net9[50] enb_bit6 avss src_out bias_pstack
x12[49] avdd pbias pcasc net9[49] enb_bit6 avss src_out bias_pstack
x12[48] avdd pbias pcasc net9[48] enb_bit6 avss src_out bias_pstack
x12[47] avdd pbias pcasc net9[47] enb_bit6 avss src_out bias_pstack
x12[46] avdd pbias pcasc net9[46] enb_bit6 avss src_out bias_pstack
x12[45] avdd pbias pcasc net9[45] enb_bit6 avss src_out bias_pstack
x12[44] avdd pbias pcasc net9[44] enb_bit6 avss src_out bias_pstack
x12[43] avdd pbias pcasc net9[43] enb_bit6 avss src_out bias_pstack
x12[42] avdd pbias pcasc net9[42] enb_bit6 avss src_out bias_pstack
x12[41] avdd pbias pcasc net9[41] enb_bit6 avss src_out bias_pstack
x12[40] avdd pbias pcasc net9[40] enb_bit6 avss src_out bias_pstack
x12[39] avdd pbias pcasc net9[39] enb_bit6 avss src_out bias_pstack
x12[38] avdd pbias pcasc net9[38] enb_bit6 avss src_out bias_pstack
x12[37] avdd pbias pcasc net9[37] enb_bit6 avss src_out bias_pstack
x12[36] avdd pbias pcasc net9[36] enb_bit6 avss src_out bias_pstack
x12[35] avdd pbias pcasc net9[35] enb_bit6 avss src_out bias_pstack
x12[34] avdd pbias pcasc net9[34] enb_bit6 avss src_out bias_pstack
x12[33] avdd pbias pcasc net9[33] enb_bit6 avss src_out bias_pstack
x12[32] avdd pbias pcasc net9[32] enb_bit6 avss src_out bias_pstack
x12[31] avdd pbias pcasc net9[31] enb_bit6 avss src_out bias_pstack
x12[30] avdd pbias pcasc net9[30] enb_bit6 avss src_out bias_pstack
x12[29] avdd pbias pcasc net9[29] enb_bit6 avss src_out bias_pstack
x12[28] avdd pbias pcasc net9[28] enb_bit6 avss src_out bias_pstack
x12[27] avdd pbias pcasc net9[27] enb_bit6 avss src_out bias_pstack
x12[26] avdd pbias pcasc net9[26] enb_bit6 avss src_out bias_pstack
x12[25] avdd pbias pcasc net9[25] enb_bit6 avss src_out bias_pstack
x12[24] avdd pbias pcasc net9[24] enb_bit6 avss src_out bias_pstack
x12[23] avdd pbias pcasc net9[23] enb_bit6 avss src_out bias_pstack
x12[22] avdd pbias pcasc net9[22] enb_bit6 avss src_out bias_pstack
x12[21] avdd pbias pcasc net9[21] enb_bit6 avss src_out bias_pstack
x12[20] avdd pbias pcasc net9[20] enb_bit6 avss src_out bias_pstack
x12[19] avdd pbias pcasc net9[19] enb_bit6 avss src_out bias_pstack
x12[18] avdd pbias pcasc net9[18] enb_bit6 avss src_out bias_pstack
x12[17] avdd pbias pcasc net9[17] enb_bit6 avss src_out bias_pstack
x12[16] avdd pbias pcasc net9[16] enb_bit6 avss src_out bias_pstack
x12[15] avdd pbias pcasc net9[15] enb_bit6 avss src_out bias_pstack
x12[14] avdd pbias pcasc net9[14] enb_bit6 avss src_out bias_pstack
x12[13] avdd pbias pcasc net9[13] enb_bit6 avss src_out bias_pstack
x12[12] avdd pbias pcasc net9[12] enb_bit6 avss src_out bias_pstack
x12[11] avdd pbias pcasc net9[11] enb_bit6 avss src_out bias_pstack
x12[10] avdd pbias pcasc net9[10] enb_bit6 avss src_out bias_pstack
x12[9] avdd pbias pcasc net9[9] enb_bit6 avss src_out bias_pstack
x12[8] avdd pbias pcasc net9[8] enb_bit6 avss src_out bias_pstack
x12[7] avdd pbias pcasc net9[7] enb_bit6 avss src_out bias_pstack
x12[6] avdd pbias pcasc net9[6] enb_bit6 avss src_out bias_pstack
x12[5] avdd pbias pcasc net9[5] enb_bit6 avss src_out bias_pstack
x12[4] avdd pbias pcasc net9[4] enb_bit6 avss src_out bias_pstack
x12[3] avdd pbias pcasc net9[3] enb_bit6 avss src_out bias_pstack
x12[2] avdd pbias pcasc net9[2] enb_bit6 avss src_out bias_pstack
x12[1] avdd pbias pcasc net9[1] enb_bit6 avss src_out bias_pstack
x12[0] avdd pbias pcasc net9[0] enb_bit6 avss src_out bias_pstack
x1[127] avdd pbias pcasc net10[127] enb_bit7 avss src_out bias_pstack
x1[126] avdd pbias pcasc net10[126] enb_bit7 avss src_out bias_pstack
x1[125] avdd pbias pcasc net10[125] enb_bit7 avss src_out bias_pstack
x1[124] avdd pbias pcasc net10[124] enb_bit7 avss src_out bias_pstack
x1[123] avdd pbias pcasc net10[123] enb_bit7 avss src_out bias_pstack
x1[122] avdd pbias pcasc net10[122] enb_bit7 avss src_out bias_pstack
x1[121] avdd pbias pcasc net10[121] enb_bit7 avss src_out bias_pstack
x1[120] avdd pbias pcasc net10[120] enb_bit7 avss src_out bias_pstack
x1[119] avdd pbias pcasc net10[119] enb_bit7 avss src_out bias_pstack
x1[118] avdd pbias pcasc net10[118] enb_bit7 avss src_out bias_pstack
x1[117] avdd pbias pcasc net10[117] enb_bit7 avss src_out bias_pstack
x1[116] avdd pbias pcasc net10[116] enb_bit7 avss src_out bias_pstack
x1[115] avdd pbias pcasc net10[115] enb_bit7 avss src_out bias_pstack
x1[114] avdd pbias pcasc net10[114] enb_bit7 avss src_out bias_pstack
x1[113] avdd pbias pcasc net10[113] enb_bit7 avss src_out bias_pstack
x1[112] avdd pbias pcasc net10[112] enb_bit7 avss src_out bias_pstack
x1[111] avdd pbias pcasc net10[111] enb_bit7 avss src_out bias_pstack
x1[110] avdd pbias pcasc net10[110] enb_bit7 avss src_out bias_pstack
x1[109] avdd pbias pcasc net10[109] enb_bit7 avss src_out bias_pstack
x1[108] avdd pbias pcasc net10[108] enb_bit7 avss src_out bias_pstack
x1[107] avdd pbias pcasc net10[107] enb_bit7 avss src_out bias_pstack
x1[106] avdd pbias pcasc net10[106] enb_bit7 avss src_out bias_pstack
x1[105] avdd pbias pcasc net10[105] enb_bit7 avss src_out bias_pstack
x1[104] avdd pbias pcasc net10[104] enb_bit7 avss src_out bias_pstack
x1[103] avdd pbias pcasc net10[103] enb_bit7 avss src_out bias_pstack
x1[102] avdd pbias pcasc net10[102] enb_bit7 avss src_out bias_pstack
x1[101] avdd pbias pcasc net10[101] enb_bit7 avss src_out bias_pstack
x1[100] avdd pbias pcasc net10[100] enb_bit7 avss src_out bias_pstack
x1[99] avdd pbias pcasc net10[99] enb_bit7 avss src_out bias_pstack
x1[98] avdd pbias pcasc net10[98] enb_bit7 avss src_out bias_pstack
x1[97] avdd pbias pcasc net10[97] enb_bit7 avss src_out bias_pstack
x1[96] avdd pbias pcasc net10[96] enb_bit7 avss src_out bias_pstack
x1[95] avdd pbias pcasc net10[95] enb_bit7 avss src_out bias_pstack
x1[94] avdd pbias pcasc net10[94] enb_bit7 avss src_out bias_pstack
x1[93] avdd pbias pcasc net10[93] enb_bit7 avss src_out bias_pstack
x1[92] avdd pbias pcasc net10[92] enb_bit7 avss src_out bias_pstack
x1[91] avdd pbias pcasc net10[91] enb_bit7 avss src_out bias_pstack
x1[90] avdd pbias pcasc net10[90] enb_bit7 avss src_out bias_pstack
x1[89] avdd pbias pcasc net10[89] enb_bit7 avss src_out bias_pstack
x1[88] avdd pbias pcasc net10[88] enb_bit7 avss src_out bias_pstack
x1[87] avdd pbias pcasc net10[87] enb_bit7 avss src_out bias_pstack
x1[86] avdd pbias pcasc net10[86] enb_bit7 avss src_out bias_pstack
x1[85] avdd pbias pcasc net10[85] enb_bit7 avss src_out bias_pstack
x1[84] avdd pbias pcasc net10[84] enb_bit7 avss src_out bias_pstack
x1[83] avdd pbias pcasc net10[83] enb_bit7 avss src_out bias_pstack
x1[82] avdd pbias pcasc net10[82] enb_bit7 avss src_out bias_pstack
x1[81] avdd pbias pcasc net10[81] enb_bit7 avss src_out bias_pstack
x1[80] avdd pbias pcasc net10[80] enb_bit7 avss src_out bias_pstack
x1[79] avdd pbias pcasc net10[79] enb_bit7 avss src_out bias_pstack
x1[78] avdd pbias pcasc net10[78] enb_bit7 avss src_out bias_pstack
x1[77] avdd pbias pcasc net10[77] enb_bit7 avss src_out bias_pstack
x1[76] avdd pbias pcasc net10[76] enb_bit7 avss src_out bias_pstack
x1[75] avdd pbias pcasc net10[75] enb_bit7 avss src_out bias_pstack
x1[74] avdd pbias pcasc net10[74] enb_bit7 avss src_out bias_pstack
x1[73] avdd pbias pcasc net10[73] enb_bit7 avss src_out bias_pstack
x1[72] avdd pbias pcasc net10[72] enb_bit7 avss src_out bias_pstack
x1[71] avdd pbias pcasc net10[71] enb_bit7 avss src_out bias_pstack
x1[70] avdd pbias pcasc net10[70] enb_bit7 avss src_out bias_pstack
x1[69] avdd pbias pcasc net10[69] enb_bit7 avss src_out bias_pstack
x1[68] avdd pbias pcasc net10[68] enb_bit7 avss src_out bias_pstack
x1[67] avdd pbias pcasc net10[67] enb_bit7 avss src_out bias_pstack
x1[66] avdd pbias pcasc net10[66] enb_bit7 avss src_out bias_pstack
x1[65] avdd pbias pcasc net10[65] enb_bit7 avss src_out bias_pstack
x1[64] avdd pbias pcasc net10[64] enb_bit7 avss src_out bias_pstack
x1[63] avdd pbias pcasc net10[63] enb_bit7 avss src_out bias_pstack
x1[62] avdd pbias pcasc net10[62] enb_bit7 avss src_out bias_pstack
x1[61] avdd pbias pcasc net10[61] enb_bit7 avss src_out bias_pstack
x1[60] avdd pbias pcasc net10[60] enb_bit7 avss src_out bias_pstack
x1[59] avdd pbias pcasc net10[59] enb_bit7 avss src_out bias_pstack
x1[58] avdd pbias pcasc net10[58] enb_bit7 avss src_out bias_pstack
x1[57] avdd pbias pcasc net10[57] enb_bit7 avss src_out bias_pstack
x1[56] avdd pbias pcasc net10[56] enb_bit7 avss src_out bias_pstack
x1[55] avdd pbias pcasc net10[55] enb_bit7 avss src_out bias_pstack
x1[54] avdd pbias pcasc net10[54] enb_bit7 avss src_out bias_pstack
x1[53] avdd pbias pcasc net10[53] enb_bit7 avss src_out bias_pstack
x1[52] avdd pbias pcasc net10[52] enb_bit7 avss src_out bias_pstack
x1[51] avdd pbias pcasc net10[51] enb_bit7 avss src_out bias_pstack
x1[50] avdd pbias pcasc net10[50] enb_bit7 avss src_out bias_pstack
x1[49] avdd pbias pcasc net10[49] enb_bit7 avss src_out bias_pstack
x1[48] avdd pbias pcasc net10[48] enb_bit7 avss src_out bias_pstack
x1[47] avdd pbias pcasc net10[47] enb_bit7 avss src_out bias_pstack
x1[46] avdd pbias pcasc net10[46] enb_bit7 avss src_out bias_pstack
x1[45] avdd pbias pcasc net10[45] enb_bit7 avss src_out bias_pstack
x1[44] avdd pbias pcasc net10[44] enb_bit7 avss src_out bias_pstack
x1[43] avdd pbias pcasc net10[43] enb_bit7 avss src_out bias_pstack
x1[42] avdd pbias pcasc net10[42] enb_bit7 avss src_out bias_pstack
x1[41] avdd pbias pcasc net10[41] enb_bit7 avss src_out bias_pstack
x1[40] avdd pbias pcasc net10[40] enb_bit7 avss src_out bias_pstack
x1[39] avdd pbias pcasc net10[39] enb_bit7 avss src_out bias_pstack
x1[38] avdd pbias pcasc net10[38] enb_bit7 avss src_out bias_pstack
x1[37] avdd pbias pcasc net10[37] enb_bit7 avss src_out bias_pstack
x1[36] avdd pbias pcasc net10[36] enb_bit7 avss src_out bias_pstack
x1[35] avdd pbias pcasc net10[35] enb_bit7 avss src_out bias_pstack
x1[34] avdd pbias pcasc net10[34] enb_bit7 avss src_out bias_pstack
x1[33] avdd pbias pcasc net10[33] enb_bit7 avss src_out bias_pstack
x1[32] avdd pbias pcasc net10[32] enb_bit7 avss src_out bias_pstack
x1[31] avdd pbias pcasc net10[31] enb_bit7 avss src_out bias_pstack
x1[30] avdd pbias pcasc net10[30] enb_bit7 avss src_out bias_pstack
x1[29] avdd pbias pcasc net10[29] enb_bit7 avss src_out bias_pstack
x1[28] avdd pbias pcasc net10[28] enb_bit7 avss src_out bias_pstack
x1[27] avdd pbias pcasc net10[27] enb_bit7 avss src_out bias_pstack
x1[26] avdd pbias pcasc net10[26] enb_bit7 avss src_out bias_pstack
x1[25] avdd pbias pcasc net10[25] enb_bit7 avss src_out bias_pstack
x1[24] avdd pbias pcasc net10[24] enb_bit7 avss src_out bias_pstack
x1[23] avdd pbias pcasc net10[23] enb_bit7 avss src_out bias_pstack
x1[22] avdd pbias pcasc net10[22] enb_bit7 avss src_out bias_pstack
x1[21] avdd pbias pcasc net10[21] enb_bit7 avss src_out bias_pstack
x1[20] avdd pbias pcasc net10[20] enb_bit7 avss src_out bias_pstack
x1[19] avdd pbias pcasc net10[19] enb_bit7 avss src_out bias_pstack
x1[18] avdd pbias pcasc net10[18] enb_bit7 avss src_out bias_pstack
x1[17] avdd pbias pcasc net10[17] enb_bit7 avss src_out bias_pstack
x1[16] avdd pbias pcasc net10[16] enb_bit7 avss src_out bias_pstack
x1[15] avdd pbias pcasc net10[15] enb_bit7 avss src_out bias_pstack
x1[14] avdd pbias pcasc net10[14] enb_bit7 avss src_out bias_pstack
x1[13] avdd pbias pcasc net10[13] enb_bit7 avss src_out bias_pstack
x1[12] avdd pbias pcasc net10[12] enb_bit7 avss src_out bias_pstack
x1[11] avdd pbias pcasc net10[11] enb_bit7 avss src_out bias_pstack
x1[10] avdd pbias pcasc net10[10] enb_bit7 avss src_out bias_pstack
x1[9] avdd pbias pcasc net10[9] enb_bit7 avss src_out bias_pstack
x1[8] avdd pbias pcasc net10[8] enb_bit7 avss src_out bias_pstack
x1[7] avdd pbias pcasc net10[7] enb_bit7 avss src_out bias_pstack
x1[6] avdd pbias pcasc net10[6] enb_bit7 avss src_out bias_pstack
x1[5] avdd pbias pcasc net10[5] enb_bit7 avss src_out bias_pstack
x1[4] avdd pbias pcasc net10[4] enb_bit7 avss src_out bias_pstack
x1[3] avdd pbias pcasc net10[3] enb_bit7 avss src_out bias_pstack
x1[2] avdd pbias pcasc net10[2] enb_bit7 avss src_out bias_pstack
x1[1] avdd pbias pcasc net10[1] enb_bit7 avss src_out bias_pstack
x1[0] avdd pbias pcasc net10[0] enb_bit7 avss src_out bias_pstack
x12 ena[0] dvdd dvss dvss avdd avdd ena_bit0 sky130_fd_sc_hvl__lsbuflv2hv_1
x14 ena[1] dvdd dvss dvss avdd avdd ena_bit1 sky130_fd_sc_hvl__lsbuflv2hv_1
x15 ena[2] dvdd dvss dvss avdd avdd ena_bit2 sky130_fd_sc_hvl__lsbuflv2hv_1
x16 ena[3] dvdd dvss dvss avdd avdd ena_bit3 sky130_fd_sc_hvl__lsbuflv2hv_1
x17 ena[4] dvdd dvss dvss avdd avdd ena_bit4 sky130_fd_sc_hvl__lsbuflv2hv_1
x18 ena[5] dvdd dvss dvss avdd avdd ena_bit5 sky130_fd_sc_hvl__lsbuflv2hv_1
x19 ena[6] dvdd dvss dvss avdd avdd ena_bit6 sky130_fd_sc_hvl__lsbuflv2hv_1
x20 ena[7] dvdd dvss dvss avdd avdd ena_bit7 sky130_fd_sc_hvl__lsbuflv2hv_1
x25 ena_bit0 dvss dvss avdd avdd enb_bit0 sky130_fd_sc_hvl__inv_2
x26 ena_bit1 dvss dvss avdd avdd enb_bit1 sky130_fd_sc_hvl__inv_2
x27 ena_bit2 dvss dvss avdd avdd enb_bit2 sky130_fd_sc_hvl__inv_2
x28 ena_bit3 dvss dvss avdd avdd enb_bit3 sky130_fd_sc_hvl__inv_2
x29 ena_bit4 dvss dvss avdd avdd enb_bit4 sky130_fd_sc_hvl__inv_2
x30 ena_bit5 dvss dvss avdd avdd enb_bit5 sky130_fd_sc_hvl__inv_2
x31 ena_bit6 dvss dvss avdd avdd enb_bit6 sky130_fd_sc_hvl__inv_2
x32 ena_bit7 dvss dvss avdd avdd enb_bit7 sky130_fd_sc_hvl__inv_2
* noconn #net2
* noconn #net1
* noconn #net3
* noconn #net4
* noconn #net5
* noconn #net6
* noconn #net7
* noconn #net8
* noconn #net9
* noconn #net10
x2 snk_out ena_bit0 net11 nbias avss bias_nstack
* noconn #net11
x2[1] snk_out ena_bit1 net12[1] nbias avss bias_nstack
x2[0] snk_out ena_bit1 net12[0] nbias avss bias_nstack
* noconn #net12
x3[3] snk_out ena_bit2 net13[3] nbias avss bias_nstack
x3[2] snk_out ena_bit2 net13[2] nbias avss bias_nstack
x3[1] snk_out ena_bit2 net13[1] nbias avss bias_nstack
x3[0] snk_out ena_bit2 net13[0] nbias avss bias_nstack
* noconn #net13
x9[7] snk_out ena_bit3 net14[7] nbias avss bias_nstack
x9[6] snk_out ena_bit3 net14[6] nbias avss bias_nstack
x9[5] snk_out ena_bit3 net14[5] nbias avss bias_nstack
x9[4] snk_out ena_bit3 net14[4] nbias avss bias_nstack
x9[3] snk_out ena_bit3 net14[3] nbias avss bias_nstack
x9[2] snk_out ena_bit3 net14[2] nbias avss bias_nstack
x9[1] snk_out ena_bit3 net14[1] nbias avss bias_nstack
x9[0] snk_out ena_bit3 net14[0] nbias avss bias_nstack
* noconn #net14
x10[15] snk_out ena_bit4 net15[15] nbias avss bias_nstack
x10[14] snk_out ena_bit4 net15[14] nbias avss bias_nstack
x10[13] snk_out ena_bit4 net15[13] nbias avss bias_nstack
x10[12] snk_out ena_bit4 net15[12] nbias avss bias_nstack
x10[11] snk_out ena_bit4 net15[11] nbias avss bias_nstack
x10[10] snk_out ena_bit4 net15[10] nbias avss bias_nstack
x10[9] snk_out ena_bit4 net15[9] nbias avss bias_nstack
x10[8] snk_out ena_bit4 net15[8] nbias avss bias_nstack
x10[7] snk_out ena_bit4 net15[7] nbias avss bias_nstack
x10[6] snk_out ena_bit4 net15[6] nbias avss bias_nstack
x10[5] snk_out ena_bit4 net15[5] nbias avss bias_nstack
x10[4] snk_out ena_bit4 net15[4] nbias avss bias_nstack
x10[3] snk_out ena_bit4 net15[3] nbias avss bias_nstack
x10[2] snk_out ena_bit4 net15[2] nbias avss bias_nstack
x10[1] snk_out ena_bit4 net15[1] nbias avss bias_nstack
x10[0] snk_out ena_bit4 net15[0] nbias avss bias_nstack
* noconn #net15
x13[31] snk_out ena_bit5 net16[31] nbias avss bias_nstack
x13[30] snk_out ena_bit5 net16[30] nbias avss bias_nstack
x13[29] snk_out ena_bit5 net16[29] nbias avss bias_nstack
x13[28] snk_out ena_bit5 net16[28] nbias avss bias_nstack
x13[27] snk_out ena_bit5 net16[27] nbias avss bias_nstack
x13[26] snk_out ena_bit5 net16[26] nbias avss bias_nstack
x13[25] snk_out ena_bit5 net16[25] nbias avss bias_nstack
x13[24] snk_out ena_bit5 net16[24] nbias avss bias_nstack
x13[23] snk_out ena_bit5 net16[23] nbias avss bias_nstack
x13[22] snk_out ena_bit5 net16[22] nbias avss bias_nstack
x13[21] snk_out ena_bit5 net16[21] nbias avss bias_nstack
x13[20] snk_out ena_bit5 net16[20] nbias avss bias_nstack
x13[19] snk_out ena_bit5 net16[19] nbias avss bias_nstack
x13[18] snk_out ena_bit5 net16[18] nbias avss bias_nstack
x13[17] snk_out ena_bit5 net16[17] nbias avss bias_nstack
x13[16] snk_out ena_bit5 net16[16] nbias avss bias_nstack
x13[15] snk_out ena_bit5 net16[15] nbias avss bias_nstack
x13[14] snk_out ena_bit5 net16[14] nbias avss bias_nstack
x13[13] snk_out ena_bit5 net16[13] nbias avss bias_nstack
x13[12] snk_out ena_bit5 net16[12] nbias avss bias_nstack
x13[11] snk_out ena_bit5 net16[11] nbias avss bias_nstack
x13[10] snk_out ena_bit5 net16[10] nbias avss bias_nstack
x13[9] snk_out ena_bit5 net16[9] nbias avss bias_nstack
x13[8] snk_out ena_bit5 net16[8] nbias avss bias_nstack
x13[7] snk_out ena_bit5 net16[7] nbias avss bias_nstack
x13[6] snk_out ena_bit5 net16[6] nbias avss bias_nstack
x13[5] snk_out ena_bit5 net16[5] nbias avss bias_nstack
x13[4] snk_out ena_bit5 net16[4] nbias avss bias_nstack
x13[3] snk_out ena_bit5 net16[3] nbias avss bias_nstack
x13[2] snk_out ena_bit5 net16[2] nbias avss bias_nstack
x13[1] snk_out ena_bit5 net16[1] nbias avss bias_nstack
x13[0] snk_out ena_bit5 net16[0] nbias avss bias_nstack
* noconn #net16
x14[63] snk_out ena_bit6 net17[63] nbias avss bias_nstack
x14[62] snk_out ena_bit6 net17[62] nbias avss bias_nstack
x14[61] snk_out ena_bit6 net17[61] nbias avss bias_nstack
x14[60] snk_out ena_bit6 net17[60] nbias avss bias_nstack
x14[59] snk_out ena_bit6 net17[59] nbias avss bias_nstack
x14[58] snk_out ena_bit6 net17[58] nbias avss bias_nstack
x14[57] snk_out ena_bit6 net17[57] nbias avss bias_nstack
x14[56] snk_out ena_bit6 net17[56] nbias avss bias_nstack
x14[55] snk_out ena_bit6 net17[55] nbias avss bias_nstack
x14[54] snk_out ena_bit6 net17[54] nbias avss bias_nstack
x14[53] snk_out ena_bit6 net17[53] nbias avss bias_nstack
x14[52] snk_out ena_bit6 net17[52] nbias avss bias_nstack
x14[51] snk_out ena_bit6 net17[51] nbias avss bias_nstack
x14[50] snk_out ena_bit6 net17[50] nbias avss bias_nstack
x14[49] snk_out ena_bit6 net17[49] nbias avss bias_nstack
x14[48] snk_out ena_bit6 net17[48] nbias avss bias_nstack
x14[47] snk_out ena_bit6 net17[47] nbias avss bias_nstack
x14[46] snk_out ena_bit6 net17[46] nbias avss bias_nstack
x14[45] snk_out ena_bit6 net17[45] nbias avss bias_nstack
x14[44] snk_out ena_bit6 net17[44] nbias avss bias_nstack
x14[43] snk_out ena_bit6 net17[43] nbias avss bias_nstack
x14[42] snk_out ena_bit6 net17[42] nbias avss bias_nstack
x14[41] snk_out ena_bit6 net17[41] nbias avss bias_nstack
x14[40] snk_out ena_bit6 net17[40] nbias avss bias_nstack
x14[39] snk_out ena_bit6 net17[39] nbias avss bias_nstack
x14[38] snk_out ena_bit6 net17[38] nbias avss bias_nstack
x14[37] snk_out ena_bit6 net17[37] nbias avss bias_nstack
x14[36] snk_out ena_bit6 net17[36] nbias avss bias_nstack
x14[35] snk_out ena_bit6 net17[35] nbias avss bias_nstack
x14[34] snk_out ena_bit6 net17[34] nbias avss bias_nstack
x14[33] snk_out ena_bit6 net17[33] nbias avss bias_nstack
x14[32] snk_out ena_bit6 net17[32] nbias avss bias_nstack
x14[31] snk_out ena_bit6 net17[31] nbias avss bias_nstack
x14[30] snk_out ena_bit6 net17[30] nbias avss bias_nstack
x14[29] snk_out ena_bit6 net17[29] nbias avss bias_nstack
x14[28] snk_out ena_bit6 net17[28] nbias avss bias_nstack
x14[27] snk_out ena_bit6 net17[27] nbias avss bias_nstack
x14[26] snk_out ena_bit6 net17[26] nbias avss bias_nstack
x14[25] snk_out ena_bit6 net17[25] nbias avss bias_nstack
x14[24] snk_out ena_bit6 net17[24] nbias avss bias_nstack
x14[23] snk_out ena_bit6 net17[23] nbias avss bias_nstack
x14[22] snk_out ena_bit6 net17[22] nbias avss bias_nstack
x14[21] snk_out ena_bit6 net17[21] nbias avss bias_nstack
x14[20] snk_out ena_bit6 net17[20] nbias avss bias_nstack
x14[19] snk_out ena_bit6 net17[19] nbias avss bias_nstack
x14[18] snk_out ena_bit6 net17[18] nbias avss bias_nstack
x14[17] snk_out ena_bit6 net17[17] nbias avss bias_nstack
x14[16] snk_out ena_bit6 net17[16] nbias avss bias_nstack
x14[15] snk_out ena_bit6 net17[15] nbias avss bias_nstack
x14[14] snk_out ena_bit6 net17[14] nbias avss bias_nstack
x14[13] snk_out ena_bit6 net17[13] nbias avss bias_nstack
x14[12] snk_out ena_bit6 net17[12] nbias avss bias_nstack
x14[11] snk_out ena_bit6 net17[11] nbias avss bias_nstack
x14[10] snk_out ena_bit6 net17[10] nbias avss bias_nstack
x14[9] snk_out ena_bit6 net17[9] nbias avss bias_nstack
x14[8] snk_out ena_bit6 net17[8] nbias avss bias_nstack
x14[7] snk_out ena_bit6 net17[7] nbias avss bias_nstack
x14[6] snk_out ena_bit6 net17[6] nbias avss bias_nstack
x14[5] snk_out ena_bit6 net17[5] nbias avss bias_nstack
x14[4] snk_out ena_bit6 net17[4] nbias avss bias_nstack
x14[3] snk_out ena_bit6 net17[3] nbias avss bias_nstack
x14[2] snk_out ena_bit6 net17[2] nbias avss bias_nstack
x14[1] snk_out ena_bit6 net17[1] nbias avss bias_nstack
x14[0] snk_out ena_bit6 net17[0] nbias avss bias_nstack
* noconn #net17
x15[127] snk_out ena_bit7 net18[127] nbias avss bias_nstack
x15[126] snk_out ena_bit7 net18[126] nbias avss bias_nstack
x15[125] snk_out ena_bit7 net18[125] nbias avss bias_nstack
x15[124] snk_out ena_bit7 net18[124] nbias avss bias_nstack
x15[123] snk_out ena_bit7 net18[123] nbias avss bias_nstack
x15[122] snk_out ena_bit7 net18[122] nbias avss bias_nstack
x15[121] snk_out ena_bit7 net18[121] nbias avss bias_nstack
x15[120] snk_out ena_bit7 net18[120] nbias avss bias_nstack
x15[119] snk_out ena_bit7 net18[119] nbias avss bias_nstack
x15[118] snk_out ena_bit7 net18[118] nbias avss bias_nstack
x15[117] snk_out ena_bit7 net18[117] nbias avss bias_nstack
x15[116] snk_out ena_bit7 net18[116] nbias avss bias_nstack
x15[115] snk_out ena_bit7 net18[115] nbias avss bias_nstack
x15[114] snk_out ena_bit7 net18[114] nbias avss bias_nstack
x15[113] snk_out ena_bit7 net18[113] nbias avss bias_nstack
x15[112] snk_out ena_bit7 net18[112] nbias avss bias_nstack
x15[111] snk_out ena_bit7 net18[111] nbias avss bias_nstack
x15[110] snk_out ena_bit7 net18[110] nbias avss bias_nstack
x15[109] snk_out ena_bit7 net18[109] nbias avss bias_nstack
x15[108] snk_out ena_bit7 net18[108] nbias avss bias_nstack
x15[107] snk_out ena_bit7 net18[107] nbias avss bias_nstack
x15[106] snk_out ena_bit7 net18[106] nbias avss bias_nstack
x15[105] snk_out ena_bit7 net18[105] nbias avss bias_nstack
x15[104] snk_out ena_bit7 net18[104] nbias avss bias_nstack
x15[103] snk_out ena_bit7 net18[103] nbias avss bias_nstack
x15[102] snk_out ena_bit7 net18[102] nbias avss bias_nstack
x15[101] snk_out ena_bit7 net18[101] nbias avss bias_nstack
x15[100] snk_out ena_bit7 net18[100] nbias avss bias_nstack
x15[99] snk_out ena_bit7 net18[99] nbias avss bias_nstack
x15[98] snk_out ena_bit7 net18[98] nbias avss bias_nstack
x15[97] snk_out ena_bit7 net18[97] nbias avss bias_nstack
x15[96] snk_out ena_bit7 net18[96] nbias avss bias_nstack
x15[95] snk_out ena_bit7 net18[95] nbias avss bias_nstack
x15[94] snk_out ena_bit7 net18[94] nbias avss bias_nstack
x15[93] snk_out ena_bit7 net18[93] nbias avss bias_nstack
x15[92] snk_out ena_bit7 net18[92] nbias avss bias_nstack
x15[91] snk_out ena_bit7 net18[91] nbias avss bias_nstack
x15[90] snk_out ena_bit7 net18[90] nbias avss bias_nstack
x15[89] snk_out ena_bit7 net18[89] nbias avss bias_nstack
x15[88] snk_out ena_bit7 net18[88] nbias avss bias_nstack
x15[87] snk_out ena_bit7 net18[87] nbias avss bias_nstack
x15[86] snk_out ena_bit7 net18[86] nbias avss bias_nstack
x15[85] snk_out ena_bit7 net18[85] nbias avss bias_nstack
x15[84] snk_out ena_bit7 net18[84] nbias avss bias_nstack
x15[83] snk_out ena_bit7 net18[83] nbias avss bias_nstack
x15[82] snk_out ena_bit7 net18[82] nbias avss bias_nstack
x15[81] snk_out ena_bit7 net18[81] nbias avss bias_nstack
x15[80] snk_out ena_bit7 net18[80] nbias avss bias_nstack
x15[79] snk_out ena_bit7 net18[79] nbias avss bias_nstack
x15[78] snk_out ena_bit7 net18[78] nbias avss bias_nstack
x15[77] snk_out ena_bit7 net18[77] nbias avss bias_nstack
x15[76] snk_out ena_bit7 net18[76] nbias avss bias_nstack
x15[75] snk_out ena_bit7 net18[75] nbias avss bias_nstack
x15[74] snk_out ena_bit7 net18[74] nbias avss bias_nstack
x15[73] snk_out ena_bit7 net18[73] nbias avss bias_nstack
x15[72] snk_out ena_bit7 net18[72] nbias avss bias_nstack
x15[71] snk_out ena_bit7 net18[71] nbias avss bias_nstack
x15[70] snk_out ena_bit7 net18[70] nbias avss bias_nstack
x15[69] snk_out ena_bit7 net18[69] nbias avss bias_nstack
x15[68] snk_out ena_bit7 net18[68] nbias avss bias_nstack
x15[67] snk_out ena_bit7 net18[67] nbias avss bias_nstack
x15[66] snk_out ena_bit7 net18[66] nbias avss bias_nstack
x15[65] snk_out ena_bit7 net18[65] nbias avss bias_nstack
x15[64] snk_out ena_bit7 net18[64] nbias avss bias_nstack
x15[63] snk_out ena_bit7 net18[63] nbias avss bias_nstack
x15[62] snk_out ena_bit7 net18[62] nbias avss bias_nstack
x15[61] snk_out ena_bit7 net18[61] nbias avss bias_nstack
x15[60] snk_out ena_bit7 net18[60] nbias avss bias_nstack
x15[59] snk_out ena_bit7 net18[59] nbias avss bias_nstack
x15[58] snk_out ena_bit7 net18[58] nbias avss bias_nstack
x15[57] snk_out ena_bit7 net18[57] nbias avss bias_nstack
x15[56] snk_out ena_bit7 net18[56] nbias avss bias_nstack
x15[55] snk_out ena_bit7 net18[55] nbias avss bias_nstack
x15[54] snk_out ena_bit7 net18[54] nbias avss bias_nstack
x15[53] snk_out ena_bit7 net18[53] nbias avss bias_nstack
x15[52] snk_out ena_bit7 net18[52] nbias avss bias_nstack
x15[51] snk_out ena_bit7 net18[51] nbias avss bias_nstack
x15[50] snk_out ena_bit7 net18[50] nbias avss bias_nstack
x15[49] snk_out ena_bit7 net18[49] nbias avss bias_nstack
x15[48] snk_out ena_bit7 net18[48] nbias avss bias_nstack
x15[47] snk_out ena_bit7 net18[47] nbias avss bias_nstack
x15[46] snk_out ena_bit7 net18[46] nbias avss bias_nstack
x15[45] snk_out ena_bit7 net18[45] nbias avss bias_nstack
x15[44] snk_out ena_bit7 net18[44] nbias avss bias_nstack
x15[43] snk_out ena_bit7 net18[43] nbias avss bias_nstack
x15[42] snk_out ena_bit7 net18[42] nbias avss bias_nstack
x15[41] snk_out ena_bit7 net18[41] nbias avss bias_nstack
x15[40] snk_out ena_bit7 net18[40] nbias avss bias_nstack
x15[39] snk_out ena_bit7 net18[39] nbias avss bias_nstack
x15[38] snk_out ena_bit7 net18[38] nbias avss bias_nstack
x15[37] snk_out ena_bit7 net18[37] nbias avss bias_nstack
x15[36] snk_out ena_bit7 net18[36] nbias avss bias_nstack
x15[35] snk_out ena_bit7 net18[35] nbias avss bias_nstack
x15[34] snk_out ena_bit7 net18[34] nbias avss bias_nstack
x15[33] snk_out ena_bit7 net18[33] nbias avss bias_nstack
x15[32] snk_out ena_bit7 net18[32] nbias avss bias_nstack
x15[31] snk_out ena_bit7 net18[31] nbias avss bias_nstack
x15[30] snk_out ena_bit7 net18[30] nbias avss bias_nstack
x15[29] snk_out ena_bit7 net18[29] nbias avss bias_nstack
x15[28] snk_out ena_bit7 net18[28] nbias avss bias_nstack
x15[27] snk_out ena_bit7 net18[27] nbias avss bias_nstack
x15[26] snk_out ena_bit7 net18[26] nbias avss bias_nstack
x15[25] snk_out ena_bit7 net18[25] nbias avss bias_nstack
x15[24] snk_out ena_bit7 net18[24] nbias avss bias_nstack
x15[23] snk_out ena_bit7 net18[23] nbias avss bias_nstack
x15[22] snk_out ena_bit7 net18[22] nbias avss bias_nstack
x15[21] snk_out ena_bit7 net18[21] nbias avss bias_nstack
x15[20] snk_out ena_bit7 net18[20] nbias avss bias_nstack
x15[19] snk_out ena_bit7 net18[19] nbias avss bias_nstack
x15[18] snk_out ena_bit7 net18[18] nbias avss bias_nstack
x15[17] snk_out ena_bit7 net18[17] nbias avss bias_nstack
x15[16] snk_out ena_bit7 net18[16] nbias avss bias_nstack
x15[15] snk_out ena_bit7 net18[15] nbias avss bias_nstack
x15[14] snk_out ena_bit7 net18[14] nbias avss bias_nstack
x15[13] snk_out ena_bit7 net18[13] nbias avss bias_nstack
x15[12] snk_out ena_bit7 net18[12] nbias avss bias_nstack
x15[11] snk_out ena_bit7 net18[11] nbias avss bias_nstack
x15[10] snk_out ena_bit7 net18[10] nbias avss bias_nstack
x15[9] snk_out ena_bit7 net18[9] nbias avss bias_nstack
x15[8] snk_out ena_bit7 net18[8] nbias avss bias_nstack
x15[7] snk_out ena_bit7 net18[7] nbias avss bias_nstack
x15[6] snk_out ena_bit7 net18[6] nbias avss bias_nstack
x15[5] snk_out ena_bit7 net18[5] nbias avss bias_nstack
x15[4] snk_out ena_bit7 net18[4] nbias avss bias_nstack
x15[3] snk_out ena_bit7 net18[3] nbias avss bias_nstack
x15[2] snk_out ena_bit7 net18[2] nbias avss bias_nstack
x15[1] snk_out ena_bit7 net18[1] nbias avss bias_nstack
x15[0] snk_out ena_bit7 net18[0] nbias avss bias_nstack
* noconn #net18
x8[7] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x8[6] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x8[5] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x8[4] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x8[3] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x8[2] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x8[1] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x8[0] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x4 ena[0] dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x5 ena[1] dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x6 ena[2] dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x7 ena[3] dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x9 ena[4] dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x10 ena[5] dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x11 ena[6] dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x13 ena[7] dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
.ends


* expanding   symbol:  brownout_ana.sym # of pins=20
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ajc_ip__brownout/xschem/brownout_ana.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ajc_ip__brownout/xschem/brownout_ana.sch
.subckt brownout_ana vin_brout otrip_decoded[7] otrip_decoded[6] otrip_decoded[5] otrip_decoded[4] otrip_decoded[3]
+ otrip_decoded[2] otrip_decoded[1] otrip_decoded[0] vin_vunder vbg_1v2 ena avdd ibg_200n itest avss dvdd isrc_sel dvss vtrip_decoded[7]
+ vtrip_decoded[6] vtrip_decoded[5] vtrip_decoded[4] vtrip_decoded[3] vtrip_decoded[2] vtrip_decoded[1] vtrip_decoded[0] dcomp brout_filt osc_ck
+ osc_ena vunder outb outb_unbuf
*.PININFO vbg_1v2:I avdd:I avss:I dvdd:I dvss:I ena:I isrc_sel:I ibg_200n:I dcomp:O itest:O osc_ena:I osc_ck:O
*+ otrip_decoded[7:0]:I vin_brout:O outb_unbuf:I outb:O vunder:O vtrip_decoded[7:0]:I vin_vunder:O brout_filt:O
xIlvls4 dcomp3v3 dvdd dvss dvss avdd avdd vl sky130_fd_sc_hvl__lsbufhv2lv_1
xIlvls0[7] otrip_decoded[7] dvdd dvss dvss avdd avdd otrip_decoded_avdd[7] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[6] otrip_decoded[6] dvdd dvss dvss avdd avdd otrip_decoded_avdd[6] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[5] otrip_decoded[5] dvdd dvss dvss avdd avdd otrip_decoded_avdd[5] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[4] otrip_decoded[4] dvdd dvss dvss avdd avdd otrip_decoded_avdd[4] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[3] otrip_decoded[3] dvdd dvss dvss avdd avdd otrip_decoded_avdd[3] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[2] otrip_decoded[2] dvdd dvss dvss avdd avdd otrip_decoded_avdd[2] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[1] otrip_decoded[1] dvdd dvss dvss avdd avdd otrip_decoded_avdd[1] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls0[0] otrip_decoded[0] dvdd dvss dvss avdd avdd otrip_decoded_avdd[0] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls1 ena dvdd dvss dvss avdd avdd ena_avdd sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls2 isrc_sel dvdd dvss dvss avdd avdd isrc_sel_avdd sky130_fd_sc_hvl__lsbuflv2hv_1
xIrsmux avdd vin_brout ena_avdd otrip_decoded_avdd[7] otrip_decoded_avdd[6] otrip_decoded_avdd[5] otrip_decoded_avdd[4]
+ otrip_decoded_avdd[3] otrip_decoded_avdd[2] otrip_decoded_avdd[1] otrip_decoded_avdd[0] vtrip_decoded_avdd[7] vtrip_decoded_avdd[6]
+ vtrip_decoded_avdd[5] vtrip_decoded_avdd[4] vtrip_decoded_avdd[3] vtrip_decoded_avdd[2] vtrip_decoded_avdd[1] vtrip_decoded_avdd[0] vin_vunder avss
+ rstring_mux
xIcomp_brout avdd ibias0 dcomp3v3 ena_avdd vin_brout vbg_1v2 avss comparator
xIbiasgen avdd ibias0 itest ibias1 ibg_200n vbg_1v2 isrc_sel_avdd ena_avdd net7 avss ibias_gen
xIosc dvdd osc_ck osc_ena dvss rc_osc
xIinv0 outb_unbuf dvss dvss dvdd dvdd net1 sky130_fd_sc_hd__inv_4
xIinv1 net1 dvss dvss dvdd dvdd outb sky130_fd_sc_hd__inv_16
xIinv3 net3 dvss dvss dvdd dvdd net2 sky130_fd_sc_hd__inv_4
xIinv4 net2 dvss dvss dvdd dvdd vunder sky130_fd_sc_hd__inv_16
xIlvls3[7] vtrip_decoded[7] dvdd dvss dvss avdd avdd vtrip_decoded_avdd[7] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls3[6] vtrip_decoded[6] dvdd dvss dvss avdd avdd vtrip_decoded_avdd[6] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls3[5] vtrip_decoded[5] dvdd dvss dvss avdd avdd vtrip_decoded_avdd[5] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls3[4] vtrip_decoded[4] dvdd dvss dvss avdd avdd vtrip_decoded_avdd[4] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls3[3] vtrip_decoded[3] dvdd dvss dvss avdd avdd vtrip_decoded_avdd[3] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls3[2] vtrip_decoded[2] dvdd dvss dvss avdd avdd vtrip_decoded_avdd[2] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls3[1] vtrip_decoded[1] dvdd dvss dvss avdd avdd vtrip_decoded_avdd[1] sky130_fd_sc_hvl__lsbuflv2hv_1
xIlvls3[0] vtrip_decoded[0] dvdd dvss dvss avdd avdd vtrip_decoded_avdd[0] sky130_fd_sc_hvl__lsbuflv2hv_1
xIcomp_vunder avdd ibias1 net4 ena_avdd vin_vunder vbg_1v2 avss comparator
xIlvls5 net4 dvdd dvss dvss avdd avdd vlu sky130_fd_sc_hvl__lsbufhv2lv_1
xIinv2 vlu dvss dvss dvdd dvdd net3 sky130_fd_sc_hd__inv_4
xIinv5 vl dvss dvss dvdd dvdd net5 sky130_fd_sc_hd__inv_4
xIinv6 net5 dvss dvss dvdd dvdd dcomp sky130_fd_sc_hd__inv_16
XC2 dcomp_filt dvss sky130_fd_pr__cap_mim_m3_2 W=30 L=30 m=6
xIschmitt dvdd dcomp_filt vsch dvss schmitt_trigger
xIinv7 vsch dvss dvss dvdd dvdd net6 sky130_fd_sc_hd__inv_4
xIinv8 net6 dvss dvss dvdd dvdd brout_filt sky130_fd_sc_hd__inv_16
XR2 dcomp_filt vl avss sky130_fd_pr__res_xhigh_po_1p41 L=700 mult=1 m=1
XQ1 avss avss net7 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
.ends


* expanding   symbol:  audiodac_drv_ls.sym # of pins=7
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_iic_ip__audiodac_lite/xschem/audiodac_drv_ls.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_iic_ip__audiodac_lite/xschem/audiodac_drv_ls.sch
.subckt audiodac_drv_ls vdd_hi out_p out_n vdd_lo in_p in_n vss_lo
*.PININFO in_p:I in_n:I out_p:O out_n:O vdd_hi:I vss_lo:I vdd_lo:I
XM6 out_p out_n vdd_hi vdd_hi sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM5 out_n out_p vdd_hi vdd_hi sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM1 casc1 in_p vss_lo vss_lo sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=10 m=1
XM2 casc2 in_n vss_lo vss_lo sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=10 m=1
XM3 out_n vdd_lo casc1 vss_lo sky130_fd_pr__nfet_05v0_nvt L=0.9 W=50 nf=5 m=1
XM4 out_p vdd_lo casc2 vss_lo sky130_fd_pr__nfet_05v0_nvt L=0.9 W=50 nf=5 m=1
.ends


* expanding   symbol:  audiodac_drv_latch.sym # of pins=4
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_iic_ip__audiodac_lite/xschem/audiodac_drv_latch.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_iic_ip__audiodac_lite/xschem/audiodac_drv_latch.sch
.subckt audiodac_drv_latch vdd_hi in_p in_n vss
*.PININFO in_p:I in_n:I vdd_hi:I vss:I
XM19 in_n in_p vdd_hi vdd_hi sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=20 nf=2 m=1
XM18 in_n in_p vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=2 m=1
XM20 in_p in_n vdd_hi vdd_hi sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=20 nf=2 m=1
XM17 in_p in_n vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=2 m=1
.ends


* expanding   symbol:  audiodac_drv_lite_half.sym # of pins=5
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_iic_ip__audiodac_lite/xschem/audiodac_drv_lite_half.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_iic_ip__audiodac_lite/xschem/audiodac_drv_lite_half.sch
.subckt audiodac_drv_lite_half vdd_hi in out vss crosscon
*.PININFO in:I out:O vdd_hi:I vss:I crosscon:B
XM10 out drv4 vdd_hi vdd_hi sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=100 nf=10 m=4
XM9 out drv4 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=100 nf=10 m=2
XM8 drv4 crosscon vdd_hi vdd_hi sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=100 nf=10 m=1
XM7 drv4 crosscon vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=50 nf=5 m=1
XM6 crosscon drv2 vdd_hi vdd_hi sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=40 nf=4 m=1
XM5 crosscon drv2 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 nf=4 m=1
XM4 drv2 drv1 vdd_hi vdd_hi sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=2 m=1
XM3 drv2 drv1 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM2 drv1 in vdd_hi vdd_hi sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM1 drv1 in vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends


* expanding   symbol:  Parallel_10B_Block2.sym # of pins=18
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/Parallel_10B_Block2.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/Parallel_10B_Block2.sch
.subckt Parallel_10B_Block2 V6 V5 V8 V9 V7 VO1 DVDD AVDD VOUT V4 V3 V2 V1 V0 VCM DVSS AVSS VBIAS
*.PININFO VOUT:B VCM:B VO1:B V5:B V6:B V7:B V8:B V9:B V0:B V1:B V2:B V3:B V4:B AVSS:B DVSS:B VBIAS:B AVDD:B DVDD:B
VI4 AVDD net25 0
.save i(vi4)
VI6 net1 net3 0
.save i(vi6)
VI7 net8 net24 0
.save i(vi7)
.save v(vout)
VI11 net26 net6 0
.save i(vi11)
VI2 net27 net5 0
.save i(vi2)
VI1 net28 net6 0
.save i(vi1)
VI3 net29 net5 0
.save i(vi3)
VICM1 net5 VCM 0
.save i(vicm1)
VICM2 net6 net1 0
.save i(vicm2)
VI5 net30 net6 0
.save i(vi5)
VI8 net31 net5 0
.save i(vi8)
VI9 net32 net6 0
.save i(vi9)
VI10 net33 net5 0
.save i(vi10)
VI12 net34 net6 0
.save i(vi12)
VI14 net35 net5 0
.save i(vi14)
VINN2 Vx1 net8 0
.save i(vinn2)
x5 V5 DVDD net34 net35 net36 net23 DVSS AVDD AVSS Universal_R_2R_Block2
x1 V6 DVDD net32 net33 net23 net22 DVSS AVDD AVSS Universal_R_2R_Block2
x2 V7 DVDD net30 net31 net22 net21 DVSS AVDD AVSS Universal_R_2R_Block2
x3 V8 DVDD net28 net29 net21 net20 DVSS AVDD AVSS Universal_R_2R_Block2
x4 V9 DVDD net26 net27 net20 net7 DVSS AVDD AVSS Universal_R_2R_Block2
VI15 AVDD net37 0
.save i(vi15)
VI16 net8 net36 0
.save i(vi16)
.save v(vx1)
VI22 AVDD net38 0
.save i(vi22)
.save v(vx32)
VICM3 VOUT net2 0
.save i(vicm3)
VI17 net39 net13 0
.save i(vi17)
VI18 net40 net12 0
.save i(vi18)
VI19 net41 net13 0
.save i(vi19)
VI20 net42 net12 0
.save i(vi20)
VICM21 net12 VCM 0
.save i(vicm21)
VICM22 net13 net1 0
.save i(vicm22)
VI23 net43 net13 0
.save i(vi23)
VI24 net44 net12 0
.save i(vi24)
VI25 net45 net13 0
.save i(vi25)
VI26 net46 net12 0
.save i(vi26)
VI27 net47 net13 0
.save i(vi27)
VI28 net48 net12 0
.save i(vi28)
x9 V0 DVDD net47 net48 net49 net16 DVSS AVDD AVSS Universal_R_2R_Block2
x10 V1 DVDD net45 net46 net16 net17 DVSS AVDD AVSS Universal_R_2R_Block2
x11 V2 DVDD net43 net44 net17 net18 DVSS AVDD AVSS Universal_R_2R_Block2
x12 V3 DVDD net41 net42 net18 net19 DVSS AVDD AVSS Universal_R_2R_Block2
x13 V4 DVDD net39 net40 net19 net14 DVSS AVDD AVSS Universal_R_2R_Block2
VI29 net15 net49 0
.save i(vi29)
VINN1 Vx32 net15 0
.save i(vinn1)
x7 net25 VOUT net1 VCM VBIAS AVSS Output_OA
x6 net37 Vx1 net9 VCM VBIAS AVSS x1_x32_OA
x8 net38 Vx32 net10 VCM VBIAS AVSS x1_x32_OA
XR11 net10 VO1 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=20 mult=1 m=1
XR12 Vx32 net10 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=640 mult=1 m=1
XR2 net9 VO1 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=40 mult=1 m=1
XR4 Vx1 net9 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=40 mult=1 m=1
XR9 net3 net24 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=1280 mult=1 m=1
XR5 net2 net3 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=1280 mult=1 m=1
XR6 net12 net11 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=20 mult=1 m=1
XR1 net11 net14 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=20 mult=1 m=1
XR3 net4 net7 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=20 mult=1 m=1
XR7 net5 net4 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=20 mult=1 m=1
.ends


* expanding   symbol:  Input_Stage_v1.sym # of pins=7
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/Input_Stage_v1.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/Input_Stage_v1.sch
.subckt Input_Stage_v1 AVDD VINP VOUT1 VINN CM AVSS VBIAS
*.PININFO VINP:B CM:B VINN:B VOUT1:B AVDD:B AVSS:B VBIAS:B
VI13 AVDD net5 0
.save i(vi13)
VI2 AVDD net6 0
.save i(vi2)
VI3 AVDD net7 0
.save i(vi3)
.save v(voneg)
.save v(vopos)
VI1 net3 net4 0
.save i(vi1)
VI4 net4 VOUT1 0
.save i(vi4)
x1 net5 VONEG VONEG VINN VBIAS AVSS Input_Stage_OA1
x2 net7 VOPOS VOPOS VINP VBIAS AVSS Input_Stage_OA1
x3 net6 net4 net2 net1 VBIAS AVSS Input_Stage_OA2
XR7 CM VINN AVSS sky130_fd_pr__res_xhigh_po_0p35 L=860 mult=1 m=1
XR5 VINP CM AVSS sky130_fd_pr__res_xhigh_po_0p35 L=860 mult=1 m=1
XR6 CM net1 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=278 mult=1 m=1
XR8 net3 net2 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=278 mult=1 m=1
XR9 net2 VONEG AVSS sky130_fd_pr__res_xhigh_po_0p35 L=34.5 mult=1 m=1
XR10 net1 VOPOS AVSS sky130_fd_pr__res_xhigh_po_0p35 L=34.5 mult=1 m=1
.ends


* expanding   symbol:  vbias_gen_pga.sym # of pins=3
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/vbias_gen_pga.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/vbias_gen_pga.sch
.subckt vbias_gen_pga VBIAS IBIAS VSS
*.PININFO VBIAS:B VSS:B IBIAS:B
.save v(vbias)
VIBIAS net1 VBIAS 0
.save i(vibias)
XM4 VBIAS VBIAS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=1
R1 IBIAS net1 sky130_fd_pr__res_generic_m1 W=1 L=0.08 m=1
.ends


* expanding   symbol:  comparator_high_gain.sym # of pins=9
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__ccomp3v/xschem/comparator_high_gain.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__ccomp3v/xschem/comparator_high_gain.sch
.subckt comparator_high_gain VDD VBN VSS VINP VOUT VINM DVDD ena3v3 DVSS
*.PININFO VINP:I VINM:I VBN:I VDD:B VSS:B VOUT:O DVDD:B ena3v3:I DVSS:B
XM3 net1 VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM19 net2 VOUTANALOG VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM20 net2 VOUTANALOG VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM21 VOUT net2 DVDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM22 VOUT net2 DVSS DVSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM1 net4 VINM net1 net1 sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=4
XM2 net3 VINP net1 net1 sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=4
XM4 net6 VINM net4 net1 sky130_fd_pr__nfet_05v0_nvt L=1 W=5 nf=1 m=10
XM5 net5 VINP net3 net1 sky130_fd_pr__nfet_05v0_nvt L=1 W=5 nf=1 m=10
XM8 VOUTANALOG ena3v3 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM9 VOUTANALOG net5 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=10 nf=2 m=2
XM10 VOUTANALOG VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=4.8 nf=1 m=2
XM11 net8 net6 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 m=2
XM12 net7 net6 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 m=2
Vmeas net8 net6 0
.save i(vmeas)
Vmeas1 net7 net5 0
.save i(vmeas1)
.ends


* expanding   symbol:  scomp_bias.sym # of pins=4
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__ccomp3v/xschem/scomp_bias.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__ccomp3v/xschem/scomp_bias.sch
.subckt scomp_bias VDD VSS VBN ena3v3
*.PININFO VBN:O VDD:B VSS:B ena3v3:I
XM3 net1 net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=20 nf=1 m=1
XM4 net3 net1 net2 VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=20 nf=1 m=1
XM5 VBN VBN net2 VDD sky130_fd_pr__pfet_g5v0d10v5 L=15 W=1 nf=1 m=1
XM1 VBN VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XM2 net1 VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XM8 net3 ena3v3 VBN VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XR2 net2 VDD VSS sky130_fd_pr__res_high_po_1p41 L=135 mult=1 m=1
.ends


* expanding   symbol:  bandgap/bandgap.sym # of pins=5
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_cw_ip/xschem/bandgap/bandgap.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_cw_ip/xschem/bandgap/bandgap.sch
.subckt bandgap vdd vbg vss bias trim[15] trim[14] trim[13] trim[12] trim[11] trim[10] trim[9] trim[8] trim[7] trim[6] trim[5]
+ trim[4] trim[3] trim[2] trim[1] trim[0]
*.PININFO vdd:B vss:B vbg:O bias:B trim[15:0]:I
XQ2 vss vss net2 sky130_fd_pr__pnp_05v5_W0p68L0p68 m=8
XQ1 vss vss vn sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XC1 gate vss sky130_fd_pr__cap_mim_m3_1 W=10 L=10 m=8
xres vbg comp vp vn vss bg_res
XR1 net1 vp vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XM1 comp gate vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=4 nf=1 m=2
XM2 vbg gate vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=4 nf=1 m=2
xtr net1 net2 trim[15] trim[14] trim[13] trim[12] trim[11] trim[10] trim[9] trim[8] trim[7] trim[6] trim[5] trim[4] trim[3]
+ trim[2] trim[1] trim[0] vss bg_trim
xamp vdd gate vp vn vss bias se_folded_cascode_p
XM3 vs1 vbg vss vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM4 gate vs1 vss vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM5 vs1 vs2 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XC2 vs2 vss sky130_fd_pr__cap_mim_m3_1 W=10 L=10 m=3
XM6 vs2 vs2 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XM7 vss vdd vs2 vs2 sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
.ends


* expanding   symbol:  bias_generator_be4.sym # of pins=51
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/bias_generator_be4.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/bias_generator_be4.sch
.subckt bias_generator_be4 dvdd dvss en_hsxo_bias en_comp_trim_n en_ov_bias avdd en_comp_bias pcasc en_hsxo_trim_n pbias
+ en_lp1_bias en_user2_trim_n en_lp2_bias en_hgbw1_bias lp1_src_100 test_src_500 lp2_src_100 en_hgbw2_bias user_src_50 idac_src_1000
+ lsxo_src_50 hsxo_src_100 comp_src_400 hgbw2_src_100 ov_src_600 user_src_150 instr1_src_100 instr2_src_100 hgbw1_src_100 en_instr1_bias
+ en_instr2_bias en_src_test en_lsxo_bias en_snk_test nbias en_user1_bias avss en_idac_bias en_user2_bias en_comp_trim_p en_hsxo_trim_p
+ en_user2_trim_p en_lp1_trim_p en_lp2_trim_p en_hgbw1_trim_p en_hgbw2_trim_p en_instr1_trim_p en_instr2_trim_p brnout_src_200 en_brnout_bias
+ bandgap_snk_250
*.PININFO avss:B avdd:B en_hsxo_trim_n:I en_instr2_bias:I hsxo_src_100:B en_instr1_bias:I en_hgbw2_bias:I ov_src_600:B
*+ en_hgbw1_bias:I comp_src_400:B en_lp2_bias:I lp1_src_100:B en_lp1_bias:I lp2_src_100:B en_comp_bias:I hgbw1_src_100:B en_ov_bias:I
*+ hgbw2_src_100:B en_hsxo_bias:I lsxo_src_50:B dvdd:B dvss:B pcasc:I pbias:I nbias:I en_comp_trim_n:I user_src_50:B instr1_src_100:B
*+ instr2_src_100:B test_src_500:B idac_src_1000:B user_src_150:B en_snk_test:I en_user2_trim_n:I en_user2_trim_p:I en_hsxo_trim_p:I en_comp_trim_p:I
*+ en_user2_bias:I en_idac_bias:I en_src_test:I en_user1_bias:I en_lsxo_bias:I en_instr2_trim_p:I en_instr1_trim_p:I en_hgbw2_trim_p:I
*+ en_hgbw1_trim_p:I en_lp2_trim_p:I en_lp1_trim_p:I brnout_src_200:B en_brnout_bias:I bandgap_snk_250:B
x18[1] net1 avss net28[1] nbias avss bias_nstack
x18[0] net1 avss net28[0] nbias avss bias_nstack
x16[17] avdd pbias pcasc net29[17] avdd avss net2 bias_pstack
x16[16] avdd pbias pcasc net29[16] avdd avss net2 bias_pstack
x16[15] avdd pbias pcasc net29[15] avdd avss net2 bias_pstack
x16[14] avdd pbias pcasc net29[14] avdd avss net2 bias_pstack
x16[13] avdd pbias pcasc net29[13] avdd avss net2 bias_pstack
x16[12] avdd pbias pcasc net29[12] avdd avss net2 bias_pstack
x16[11] avdd pbias pcasc net29[11] avdd avss net2 bias_pstack
x16[10] avdd pbias pcasc net29[10] avdd avss net2 bias_pstack
x16[9] avdd pbias pcasc net29[9] avdd avss net2 bias_pstack
x16[8] avdd pbias pcasc net29[8] avdd avss net2 bias_pstack
x16[7] avdd pbias pcasc net29[7] avdd avss net2 bias_pstack
x16[6] avdd pbias pcasc net29[6] avdd avss net2 bias_pstack
x16[5] avdd pbias pcasc net29[5] avdd avss net2 bias_pstack
x16[4] avdd pbias pcasc net29[4] avdd avss net2 bias_pstack
x16[3] avdd pbias pcasc net29[3] avdd avss net2 bias_pstack
x16[2] avdd pbias pcasc net29[2] avdd avss net2 bias_pstack
x16[1] avdd pbias pcasc net29[1] avdd avss net2 bias_pstack
x16[0] avdd pbias pcasc net29[0] avdd avss net2 bias_pstack
x8[1] avdd pbias pcasc net30[1] enb_hsxo_3v3 avss hsxo_src_100 bias_pstack
x8[0] avdd pbias pcasc net30[0] enb_hsxo_3v3 avss hsxo_src_100 bias_pstack
x4[11] avdd pbias pcasc net31[11] enb_ov_3v3 avss ov_src_600 bias_pstack
x4[10] avdd pbias pcasc net31[10] enb_ov_3v3 avss ov_src_600 bias_pstack
x4[9] avdd pbias pcasc net31[9] enb_ov_3v3 avss ov_src_600 bias_pstack
x4[8] avdd pbias pcasc net31[8] enb_ov_3v3 avss ov_src_600 bias_pstack
x4[7] avdd pbias pcasc net31[7] enb_ov_3v3 avss ov_src_600 bias_pstack
x4[6] avdd pbias pcasc net31[6] enb_ov_3v3 avss ov_src_600 bias_pstack
x4[5] avdd pbias pcasc net31[5] enb_ov_3v3 avss ov_src_600 bias_pstack
x4[4] avdd pbias pcasc net31[4] enb_ov_3v3 avss ov_src_600 bias_pstack
x4[3] avdd pbias pcasc net31[3] enb_ov_3v3 avss ov_src_600 bias_pstack
x4[2] avdd pbias pcasc net31[2] enb_ov_3v3 avss ov_src_600 bias_pstack
x4[1] avdd pbias pcasc net31[1] enb_ov_3v3 avss ov_src_600 bias_pstack
x4[0] avdd pbias pcasc net31[0] enb_ov_3v3 avss ov_src_600 bias_pstack
x5[7] avdd pbias pcasc net32[7] enb_comp_3v3 avss comp_src_400 bias_pstack
x5[6] avdd pbias pcasc net32[6] enb_comp_3v3 avss comp_src_400 bias_pstack
x5[5] avdd pbias pcasc net32[5] enb_comp_3v3 avss comp_src_400 bias_pstack
x5[4] avdd pbias pcasc net32[4] enb_comp_3v3 avss comp_src_400 bias_pstack
x5[3] avdd pbias pcasc net32[3] enb_comp_3v3 avss comp_src_400 bias_pstack
x5[2] avdd pbias pcasc net32[2] enb_comp_3v3 avss comp_src_400 bias_pstack
x5[1] avdd pbias pcasc net32[1] enb_comp_3v3 avss comp_src_400 bias_pstack
x5[0] avdd pbias pcasc net32[0] enb_comp_3v3 avss comp_src_400 bias_pstack
x6[1] avdd pbias pcasc net33[1] enb_lp1_3v3 avss lp1_src_100 bias_pstack
x6[0] avdd pbias pcasc net33[0] enb_lp1_3v3 avss lp1_src_100 bias_pstack
x7[1] avdd pbias pcasc net34[1] enb_lp2_3v3 avss lp2_src_100 bias_pstack
x7[0] avdd pbias pcasc net34[0] enb_lp2_3v3 avss lp2_src_100 bias_pstack
x11[1] avdd pbias pcasc net35[1] enb_hgbw1_3v3 avss hgbw1_src_100 bias_pstack
x11[0] avdd pbias pcasc net35[0] enb_hgbw1_3v3 avss hgbw1_src_100 bias_pstack
x12[1] avdd pbias pcasc net36[1] enb_hgbw2_3v3 avss hgbw2_src_100 bias_pstack
x12[0] avdd pbias pcasc net36[0] enb_hgbw2_3v3 avss hgbw2_src_100 bias_pstack
x13 avdd pbias pcasc net37 enb_lsxo_3v3 avss lsxo_src_50 bias_pstack
x10 en_hsxo_trim_n dvdd dvss dvss avdd avdd ena_hsxo_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x12 en_hsxo_bias dvdd dvss dvss avdd avdd net11 sky130_fd_sc_hvl__lsbuflv2hv_1
x14 en_ov_bias dvdd dvss dvss avdd avdd net10 sky130_fd_sc_hvl__lsbuflv2hv_1
x15 en_comp_bias dvdd dvss dvss avdd avdd net9 sky130_fd_sc_hvl__lsbuflv2hv_1
x16 en_lp1_bias dvdd dvss dvss avdd avdd net8 sky130_fd_sc_hvl__lsbuflv2hv_1
x17 en_lp2_bias dvdd dvss dvss avdd avdd net7 sky130_fd_sc_hvl__lsbuflv2hv_1
x18 en_hgbw1_bias dvdd dvss dvss avdd avdd net6 sky130_fd_sc_hvl__lsbuflv2hv_1
x19 en_hgbw2_bias dvdd dvss dvss avdd avdd net5 sky130_fd_sc_hvl__lsbuflv2hv_1
x20 en_instr1_bias dvdd dvss dvss avdd avdd net4 sky130_fd_sc_hvl__lsbuflv2hv_1
x22 en_instr2_bias dvdd dvss dvss avdd avdd net3 sky130_fd_sc_hvl__lsbuflv2hv_1
x25 net11 dvss dvss avdd avdd enb_hsxo_3v3 sky130_fd_sc_hvl__inv_2
x26 net10 dvss dvss avdd avdd enb_ov_3v3 sky130_fd_sc_hvl__inv_2
x27 net9 dvss dvss avdd avdd enb_comp_3v3 sky130_fd_sc_hvl__inv_2
x28 net8 dvss dvss avdd avdd enb_lp1_3v3 sky130_fd_sc_hvl__inv_2
x29 net7 dvss dvss avdd avdd enb_lp2_3v3 sky130_fd_sc_hvl__inv_2
x30 net6 dvss dvss avdd avdd enb_hgbw1_3v3 sky130_fd_sc_hvl__inv_2
x31 net5 dvss dvss avdd avdd enb_hgbw2_3v3 sky130_fd_sc_hvl__inv_2
x32 net4 dvss dvss avdd avdd enb_instr1_3v3 sky130_fd_sc_hvl__inv_2
x34 net3 dvss dvss avdd avdd enb_instr2_3v3 sky130_fd_sc_hvl__inv_2
* noconn #net29
* noconn #net28
* noconn #net30
* noconn #net31
* noconn #net32
* noconn #net33
* noconn #net34
* noconn #net35
* noconn #net36
* noconn #net37
x1[1] comp_src_400 ena_comp_3v3 net38[1] nbias avss bias_nstack
x1[0] comp_src_400 ena_comp_3v3 net38[0] nbias avss bias_nstack
* noconn #net38
x1 en_comp_trim_n dvdd dvss dvss avdd avdd ena_comp_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x2 avdd pbias pcasc net39 enb_user1_3v3 avss user_src_50 bias_pstack
* noconn #net39
x3[1] avdd pbias pcasc net40[1] enb_instr1_3v3 avss instr1_src_100 bias_pstack
x3[0] avdd pbias pcasc net40[0] enb_instr1_3v3 avss instr1_src_100 bias_pstack
* noconn #net40
x2[1] avdd pbias pcasc net41[1] enb_instr2_3v3 avss instr2_src_100 bias_pstack
x2[0] avdd pbias pcasc net41[0] enb_instr2_3v3 avss instr2_src_100 bias_pstack
* noconn #net41
x9[9] avdd pbias pcasc net42[9] enb_test_3v3 avss test_src_500 bias_pstack
x9[8] avdd pbias pcasc net42[8] enb_test_3v3 avss test_src_500 bias_pstack
x9[7] avdd pbias pcasc net42[7] enb_test_3v3 avss test_src_500 bias_pstack
x9[6] avdd pbias pcasc net42[6] enb_test_3v3 avss test_src_500 bias_pstack
x9[5] avdd pbias pcasc net42[5] enb_test_3v3 avss test_src_500 bias_pstack
x9[4] avdd pbias pcasc net42[4] enb_test_3v3 avss test_src_500 bias_pstack
x9[3] avdd pbias pcasc net42[3] enb_test_3v3 avss test_src_500 bias_pstack
x9[2] avdd pbias pcasc net42[2] enb_test_3v3 avss test_src_500 bias_pstack
x9[1] avdd pbias pcasc net42[1] enb_test_3v3 avss test_src_500 bias_pstack
x9[0] avdd pbias pcasc net42[0] enb_test_3v3 avss test_src_500 bias_pstack
* noconn #net42
x10[19] avdd pbias pcasc net43[19] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[18] avdd pbias pcasc net43[18] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[17] avdd pbias pcasc net43[17] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[16] avdd pbias pcasc net43[16] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[15] avdd pbias pcasc net43[15] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[14] avdd pbias pcasc net43[14] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[13] avdd pbias pcasc net43[13] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[12] avdd pbias pcasc net43[12] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[11] avdd pbias pcasc net43[11] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[10] avdd pbias pcasc net43[10] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[9] avdd pbias pcasc net43[9] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[8] avdd pbias pcasc net43[8] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[7] avdd pbias pcasc net43[7] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[6] avdd pbias pcasc net43[6] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[5] avdd pbias pcasc net43[5] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[4] avdd pbias pcasc net43[4] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[3] avdd pbias pcasc net43[3] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[2] avdd pbias pcasc net43[2] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[1] avdd pbias pcasc net43[1] enb_idac_3v3 avss idac_src_1000 bias_pstack
x10[0] avdd pbias pcasc net43[0] enb_idac_3v3 avss idac_src_1000 bias_pstack
* noconn #net43
x13[1] hsxo_src_100 ena_hsxo_3v3 net44[1] nbias avss bias_nstack
x13[0] hsxo_src_100 ena_hsxo_3v3 net44[0] nbias avss bias_nstack
* noconn #net44
x14[1] user_src_150 ena_user2_3v3 net45[1] nbias avss bias_nstack
x14[0] user_src_150 ena_user2_3v3 net45[0] nbias avss bias_nstack
* noconn #net45
x15[74] test_src_500 ena_test_3v3 net46[74] nbias avss bias_nstack
x15[73] test_src_500 ena_test_3v3 net46[73] nbias avss bias_nstack
x15[72] test_src_500 ena_test_3v3 net46[72] nbias avss bias_nstack
x15[71] test_src_500 ena_test_3v3 net46[71] nbias avss bias_nstack
x15[70] test_src_500 ena_test_3v3 net46[70] nbias avss bias_nstack
x15[69] test_src_500 ena_test_3v3 net46[69] nbias avss bias_nstack
x15[68] test_src_500 ena_test_3v3 net46[68] nbias avss bias_nstack
x15[67] test_src_500 ena_test_3v3 net46[67] nbias avss bias_nstack
x15[66] test_src_500 ena_test_3v3 net46[66] nbias avss bias_nstack
x15[65] test_src_500 ena_test_3v3 net46[65] nbias avss bias_nstack
x15[64] test_src_500 ena_test_3v3 net46[64] nbias avss bias_nstack
x15[63] test_src_500 ena_test_3v3 net46[63] nbias avss bias_nstack
x15[62] test_src_500 ena_test_3v3 net46[62] nbias avss bias_nstack
x15[61] test_src_500 ena_test_3v3 net46[61] nbias avss bias_nstack
x15[60] test_src_500 ena_test_3v3 net46[60] nbias avss bias_nstack
x15[59] test_src_500 ena_test_3v3 net46[59] nbias avss bias_nstack
x15[58] test_src_500 ena_test_3v3 net46[58] nbias avss bias_nstack
x15[57] test_src_500 ena_test_3v3 net46[57] nbias avss bias_nstack
x15[56] test_src_500 ena_test_3v3 net46[56] nbias avss bias_nstack
x15[55] test_src_500 ena_test_3v3 net46[55] nbias avss bias_nstack
x15[54] test_src_500 ena_test_3v3 net46[54] nbias avss bias_nstack
x15[53] test_src_500 ena_test_3v3 net46[53] nbias avss bias_nstack
x15[52] test_src_500 ena_test_3v3 net46[52] nbias avss bias_nstack
x15[51] test_src_500 ena_test_3v3 net46[51] nbias avss bias_nstack
x15[50] test_src_500 ena_test_3v3 net46[50] nbias avss bias_nstack
x15[49] test_src_500 ena_test_3v3 net46[49] nbias avss bias_nstack
x15[48] test_src_500 ena_test_3v3 net46[48] nbias avss bias_nstack
x15[47] test_src_500 ena_test_3v3 net46[47] nbias avss bias_nstack
x15[46] test_src_500 ena_test_3v3 net46[46] nbias avss bias_nstack
x15[45] test_src_500 ena_test_3v3 net46[45] nbias avss bias_nstack
x15[44] test_src_500 ena_test_3v3 net46[44] nbias avss bias_nstack
x15[43] test_src_500 ena_test_3v3 net46[43] nbias avss bias_nstack
x15[42] test_src_500 ena_test_3v3 net46[42] nbias avss bias_nstack
x15[41] test_src_500 ena_test_3v3 net46[41] nbias avss bias_nstack
x15[40] test_src_500 ena_test_3v3 net46[40] nbias avss bias_nstack
x15[39] test_src_500 ena_test_3v3 net46[39] nbias avss bias_nstack
x15[38] test_src_500 ena_test_3v3 net46[38] nbias avss bias_nstack
x15[37] test_src_500 ena_test_3v3 net46[37] nbias avss bias_nstack
x15[36] test_src_500 ena_test_3v3 net46[36] nbias avss bias_nstack
x15[35] test_src_500 ena_test_3v3 net46[35] nbias avss bias_nstack
x15[34] test_src_500 ena_test_3v3 net46[34] nbias avss bias_nstack
x15[33] test_src_500 ena_test_3v3 net46[33] nbias avss bias_nstack
x15[32] test_src_500 ena_test_3v3 net46[32] nbias avss bias_nstack
x15[31] test_src_500 ena_test_3v3 net46[31] nbias avss bias_nstack
x15[30] test_src_500 ena_test_3v3 net46[30] nbias avss bias_nstack
x15[29] test_src_500 ena_test_3v3 net46[29] nbias avss bias_nstack
x15[28] test_src_500 ena_test_3v3 net46[28] nbias avss bias_nstack
x15[27] test_src_500 ena_test_3v3 net46[27] nbias avss bias_nstack
x15[26] test_src_500 ena_test_3v3 net46[26] nbias avss bias_nstack
x15[25] test_src_500 ena_test_3v3 net46[25] nbias avss bias_nstack
x15[24] test_src_500 ena_test_3v3 net46[24] nbias avss bias_nstack
x15[23] test_src_500 ena_test_3v3 net46[23] nbias avss bias_nstack
x15[22] test_src_500 ena_test_3v3 net46[22] nbias avss bias_nstack
x15[21] test_src_500 ena_test_3v3 net46[21] nbias avss bias_nstack
x15[20] test_src_500 ena_test_3v3 net46[20] nbias avss bias_nstack
x15[19] test_src_500 ena_test_3v3 net46[19] nbias avss bias_nstack
x15[18] test_src_500 ena_test_3v3 net46[18] nbias avss bias_nstack
x15[17] test_src_500 ena_test_3v3 net46[17] nbias avss bias_nstack
x15[16] test_src_500 ena_test_3v3 net46[16] nbias avss bias_nstack
x15[15] test_src_500 ena_test_3v3 net46[15] nbias avss bias_nstack
x15[14] test_src_500 ena_test_3v3 net46[14] nbias avss bias_nstack
x15[13] test_src_500 ena_test_3v3 net46[13] nbias avss bias_nstack
x15[12] test_src_500 ena_test_3v3 net46[12] nbias avss bias_nstack
x15[11] test_src_500 ena_test_3v3 net46[11] nbias avss bias_nstack
x15[10] test_src_500 ena_test_3v3 net46[10] nbias avss bias_nstack
x15[9] test_src_500 ena_test_3v3 net46[9] nbias avss bias_nstack
x15[8] test_src_500 ena_test_3v3 net46[8] nbias avss bias_nstack
x15[7] test_src_500 ena_test_3v3 net46[7] nbias avss bias_nstack
x15[6] test_src_500 ena_test_3v3 net46[6] nbias avss bias_nstack
x15[5] test_src_500 ena_test_3v3 net46[5] nbias avss bias_nstack
x15[4] test_src_500 ena_test_3v3 net46[4] nbias avss bias_nstack
x15[3] test_src_500 ena_test_3v3 net46[3] nbias avss bias_nstack
x15[2] test_src_500 ena_test_3v3 net46[2] nbias avss bias_nstack
x15[1] test_src_500 ena_test_3v3 net46[1] nbias avss bias_nstack
x15[0] test_src_500 ena_test_3v3 net46[0] nbias avss bias_nstack
* noconn #net46
x17[2] avdd pbias pcasc net47[2] enb_user2_3v3 avss user_src_150 bias_pstack
x17[1] avdd pbias pcasc net47[1] enb_user2_3v3 avss user_src_150 bias_pstack
x17[0] avdd pbias pcasc net47[0] enb_user2_3v3 avss user_src_150 bias_pstack
* noconn #net47
* noconn #net2
* noconn #net1
x3 avdd pbias pcasc net48 enb_comp_trim_3v3 avss comp_src_400 bias_pstack
* noconn #net48
x4 avdd pbias pcasc net49 enb_hsxo_trim_3v3 avss hsxo_src_100 bias_pstack
* noconn #net49
x5 avdd pbias pcasc net50 enb_user2_trim_3v3 avss user_src_150 bias_pstack
* noconn #net50
x6 avdd pbias pcasc net51 enb_lp1_trim_3v3 avss lp1_src_100 bias_pstack
* noconn #net51
x7 avdd pbias pcasc net52 enb_lp2_trim_3v3 avss lp2_src_100 bias_pstack
* noconn #net52
x8 avdd pbias pcasc net53 enb_hgbw1_trim_3v3 avss hgbw1_src_100 bias_pstack
* noconn #net53
x9 avdd pbias pcasc net54 enb_hgbw2_trim_3v3 avss hgbw2_src_100 bias_pstack
* noconn #net54
x11 avdd pbias pcasc net55 enb_instr1_trim_3v3 avss instr1_src_100 bias_pstack
* noconn #net55
x21 avdd pbias pcasc net56 enb_instr2_trim_3v3 avss instr2_src_100 bias_pstack
* noconn #net56
x24 en_snk_test dvdd dvss dvss avdd avdd ena_test_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x33 en_user2_trim_n dvdd dvss dvss avdd avdd ena_user2_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x35 en_lsxo_bias dvdd dvss dvss avdd avdd net18 sky130_fd_sc_hvl__lsbuflv2hv_1
x36 en_user1_bias dvdd dvss dvss avdd avdd net17 sky130_fd_sc_hvl__lsbuflv2hv_1
x37 en_src_test dvdd dvss dvss avdd avdd ena_bandgap_3v3 sky130_fd_sc_hvl__lsbuflv2hv_1
x38 en_idac_bias dvdd dvss dvss avdd avdd net16 sky130_fd_sc_hvl__lsbuflv2hv_1
x39 en_user2_bias dvdd dvss dvss avdd avdd net15 sky130_fd_sc_hvl__lsbuflv2hv_1
x40 en_comp_trim_p dvdd dvss dvss avdd avdd net14 sky130_fd_sc_hvl__lsbuflv2hv_1
x41 en_hsxo_trim_p dvdd dvss dvss avdd avdd net13 sky130_fd_sc_hvl__lsbuflv2hv_1
x42 en_user2_trim_p dvdd dvss dvss avdd avdd net12 sky130_fd_sc_hvl__lsbuflv2hv_1
x44 net18 dvss dvss avdd avdd enb_lsxo_3v3 sky130_fd_sc_hvl__inv_2
x45 net17 dvss dvss avdd avdd enb_user1_3v3 sky130_fd_sc_hvl__inv_2
x46 ena_bandgap_3v3 dvss dvss avdd avdd enb_test_3v3 sky130_fd_sc_hvl__inv_2
x47 net16 dvss dvss avdd avdd enb_idac_3v3 sky130_fd_sc_hvl__inv_2
x48 net15 dvss dvss avdd avdd enb_user2_3v3 sky130_fd_sc_hvl__inv_2
x49 net14 dvss dvss avdd avdd enb_comp_trim_3v3 sky130_fd_sc_hvl__inv_2
x50 net13 dvss dvss avdd avdd enb_hsxo_trim_3v3 sky130_fd_sc_hvl__inv_2
x51 net12 dvss dvss avdd avdd enb_user2_trim_3v3 sky130_fd_sc_hvl__inv_2
x53 en_lp1_trim_p dvdd dvss dvss avdd avdd net24 sky130_fd_sc_hvl__lsbuflv2hv_1
x54 en_lp2_trim_p dvdd dvss dvss avdd avdd net23 sky130_fd_sc_hvl__lsbuflv2hv_1
x55 en_hgbw1_trim_p dvdd dvss dvss avdd avdd net22 sky130_fd_sc_hvl__lsbuflv2hv_1
x56 en_hgbw2_trim_p dvdd dvss dvss avdd avdd net21 sky130_fd_sc_hvl__lsbuflv2hv_1
x57 en_instr1_trim_p dvdd dvss dvss avdd avdd net20 sky130_fd_sc_hvl__lsbuflv2hv_1
x58 en_instr2_trim_p dvdd dvss dvss avdd avdd net19 sky130_fd_sc_hvl__lsbuflv2hv_1
x59 net24 dvss dvss avdd avdd enb_lp1_trim_3v3 sky130_fd_sc_hvl__inv_2
x60 net23 dvss dvss avdd avdd enb_lp2_trim_3v3 sky130_fd_sc_hvl__inv_2
x61 net22 dvss dvss avdd avdd enb_hgbw1_trim_3v3 sky130_fd_sc_hvl__inv_2
x62 net21 dvss dvss avdd avdd enb_hgbw2_trim_3v3 sky130_fd_sc_hvl__inv_2
x63 net20 dvss dvss avdd avdd enb_instr1_trim_3v3 sky130_fd_sc_hvl__inv_2
x64 net19 dvss dvss avdd avdd enb_instr2_trim_3v3 sky130_fd_sc_hvl__inv_2
x19[3] avdd pbias pcasc net57[3] enb_brnout_3v3 avss brnout_src_200 bias_pstack
x19[2] avdd pbias pcasc net57[2] enb_brnout_3v3 avss brnout_src_200 bias_pstack
x19[1] avdd pbias pcasc net57[1] enb_brnout_3v3 avss brnout_src_200 bias_pstack
x19[0] avdd pbias pcasc net57[0] enb_brnout_3v3 avss brnout_src_200 bias_pstack
* noconn #net57
x65 en_brnout_bias dvdd dvss dvss avdd avdd net25 sky130_fd_sc_hvl__lsbuflv2hv_1
x66 net25 dvss dvss avdd avdd enb_brnout_3v3 sky130_fd_sc_hvl__inv_2
x23[3] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x23[2] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x23[1] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x23[0] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x20[13] net26 avss net58[13] nbias avss bias_nstack
x20[12] net26 avss net58[12] nbias avss bias_nstack
x20[11] net26 avss net58[11] nbias avss bias_nstack
x20[10] net26 avss net58[10] nbias avss bias_nstack
x20[9] net26 avss net58[9] nbias avss bias_nstack
x20[8] net26 avss net58[8] nbias avss bias_nstack
x20[7] net26 avss net58[7] nbias avss bias_nstack
x20[6] net26 avss net58[6] nbias avss bias_nstack
x20[5] net26 avss net58[5] nbias avss bias_nstack
x20[4] net26 avss net58[4] nbias avss bias_nstack
x20[3] net26 avss net58[3] nbias avss bias_nstack
x20[2] net26 avss net58[2] nbias avss bias_nstack
x20[1] net26 avss net58[1] nbias avss bias_nstack
x20[0] net26 avss net58[0] nbias avss bias_nstack
* noconn #net58
* noconn #net26
x23 en_hsxo_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x43 en_ov_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x52 en_comp_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x67 en_lp1_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x68 en_lp2_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x69 en_hgbw1_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x70 en_hgbw2_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x71 en_instr1_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x72 en_instr2_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x73 en_lsxo_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x74 en_user1_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x75 en_idac_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x76 en_user2_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x77 en_brnout_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x78 en_comp_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x79 en_hsxo_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x80 en_user2_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x81 en_lp1_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x82 en_lp2_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x83 en_hgbw1_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x84 en_hgbw2_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x85 en_instr1_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x86 en_instr2_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x87 en_comp_trim_n dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x88 en_hsxo_trim_n dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x89 en_user2_trim_n dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x90 en_src_test dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x91 en_snk_test dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
x21[4] bandgap_snk_250 ena_bandgap_3v3 net59[4] nbias avss bias_nstack
x21[3] bandgap_snk_250 ena_bandgap_3v3 net59[3] nbias avss bias_nstack
x21[2] bandgap_snk_250 ena_bandgap_3v3 net59[2] nbias avss bias_nstack
x21[1] bandgap_snk_250 ena_bandgap_3v3 net59[1] nbias avss bias_nstack
x21[0] bandgap_snk_250 ena_bandgap_3v3 net59[0] nbias avss bias_nstack
* noconn #net59
x22[1] avdd pbias pcasc net60[1] avdd avss net27 bias_pstack
x22[0] avdd pbias pcasc net60[0] avdd avss net27 bias_pstack
* noconn #net60
* noconn #net27
.ends


* expanding   symbol:  comparator_final.sym # of pins=8
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_sw_ip__por/xschem/comparator_final.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_sw_ip__por/xschem/comparator_final.sch
.subckt comparator_final Vinn Vinp RST VSS AVDD DVDD vo ibn180n
*.PININFO AVDD:I RST:O VSS:I Vinn:I Vinp:I DVDD:I vo:O ibn180n:O
XM1 VS vbn VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM3 vbp vbp AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM2 vt vbp AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM7 vo vt AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM6 vo vbn VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM14 vo1 vo VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM15 vo1 vo net1 net1 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM12 net4 vo1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM13 net4 vo1 DVDD DVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM16 RST net4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM17 RST net4 DVDD DVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM4 vbp AVDD net3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM8 vt AVDD net2 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM19 net1 net1 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM23 net5 net5 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 m=1
XM24 vbn net5 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 m=1
XR12 VSS net6 VSS sky130_fd_pr__res_xhigh_po_0p35 L=28 mult=1 m=1
XM25 vbn vbn VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM26 net5 vbn net6 VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=2
XM28 net7 vbn VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=4 nf=1 m=1
XM18 net2 Vinn VS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 m=7
XM10 net3 Vinp VS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 m=2
XM5 net8 net8 AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 m=1
XM11 net9 net9 net8 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 m=1
XM20 net7 net7 net9 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=1 nf=1 m=1
XM21 net5 net7 vbn VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM9 net10 vbn VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
Vbn180n ibn180n net10 0
.save i(vbn180n)
XM22 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=2 nf=1 m=1
.ends


* expanding   symbol:  delayPulse_final.sym # of pins=8
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_sw_ip__por/xschem/delayPulse_final.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_sw_ip__por/xschem/delayPulse_final.sch
.subckt delayPulse_final din por VCCL VSS VCCH porb porb_h[1] porb_h[0] ibn180n
*.PININFO VCCL:I VSS:I din:I por:O VCCH:I porb:O porb_h[1:0]:O ibn180n:I
x1 Td_L Td_Sd VSS VSS VCCL VCCL outxor sky130_fd_sc_ls__xor2_1
x3 porbPre porbhPre VCCL VSS VCCH levelShifter
XM2 net1 din VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 m=2
XM3 Td_S net1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 m=2
XM5 VT2 net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=2 m=1
XM7 net1 din VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=0.5 nf=1 m=2
XM8 Td_S net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=0.5 nf=1 m=2
XM10 VT2 net1 net10 VCCL sky130_fd_pr__pfet_01v8 L=0.3 W=2 nf=2 m=1
XM13 net4 VT3 VSS VSS sky130_fd_pr__nfet_01v8 L=0.3 W=0.5 nf=1 m=2
XM14 net4 VT3 net5 net5 sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 m=2
x4 net2 VSS VCCL TieH_1p8
XM11 vbn1 net8 net6 VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=2 nf=1 m=1
XM17 vbp1 vbn1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=2 nf=1 m=1
XM18 net6 net7 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=2 nf=1 m=1
XM19 vbn1 vbn1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=2 nf=1 m=7
XM24 net8 net8 net7 VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=2 nf=1 m=1
XM25 net7 net7 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=16 nf=8 m=1
XM26 VSS VSS net9 VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XM6 VT3 VT2 net3 VSS sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=2 m=1
XM12 VT3 VT2 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.3 W=2 nf=2 m=1
XM1 vbp1 vbp1 vbp1 VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 m=1
XM15 vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 m=7
XM16 net10 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 m=1
XM20 net10 vbp1 net10 VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 m=1
XM21 net3 vbn1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=2 nf=1 m=4
XM22 net5 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 m=4
XM23 net5 vbp1 net5 VCCL sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=2 m=1
XM27 net11 net4 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM29 net11 net4 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
XM30 Td_L net11 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=2
XM31 Td_L net11 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=2
XM32 net12 Td_S VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM33 net12 Td_S VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
XM34 net13 net12 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM35 net13 net12 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
XM36 Td_Sd net14 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=2
XM38 net14 net13 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM39 net14 net13 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
x6 outxor VSS VSS VCCL VCCL rstn sky130_fd_sc_ls__buf_8
XC4 VSS net13 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 m=1
XC7 VSS VT2 sky130_fd_pr__cap_mim_m3_2 W=16 L=16 m=20
XC2 VCCL VT3 sky130_fd_pr__cap_mim_m3_2 W=16 L=16 m=20
XC8 VCCL net12 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 m=1
XC9 VCCL net14 sky130_fd_pr__cap_mim_m3_2 W=10 L=10 m=1
XM40 Td_Sd net14 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=2
x5 rstn net2 Td_Sd VSS VSS VCCL VCCL porbPre sky130_fd_sc_ls__dfrtn_1
x2 Td_Sd net2 Td_Lb VSS VSS VCCL VCCL porPre sky130_fd_sc_ls__dfrtp_1
XM4 Td_Lb Td_L VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=2
XM9 Td_Lb Td_L VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=2
XC1 VSS vbn1 sky130_fd_pr__cap_mim_m3_2 W=16 L=16 m=1
XC5 VCCH net7 sky130_fd_pr__cap_mim_m3_2 W=16 L=16 m=1
XC6 VCCL vbp1 sky130_fd_pr__cap_mim_m3_2 W=16 L=16 m=1
XC3 VCCH net8 sky130_fd_pr__cap_mim_m3_2 W=8 L=8 m=1
XM28 net15 porPre VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM37 net15 porPre VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
XM41 net16 net15 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=2
XM42 net16 net15 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=2
XM43 net17 net16 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=8
XM44 net17 net16 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=8
XM45 por net17 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=16
XM46 por net17 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=16
XM47 net18 porbPre VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM48 net18 porbPre VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
XM49 net19 net18 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=2
XM50 net19 net18 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=2
XM51 net20 net19 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=8
XM52 net20 net19 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=8
XM53 porb net20 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=16
XM54 porb net20 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=16
XM59 net21 porbhPre VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM60 net21 porbhPre VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=2 m=1
x7 VSS VSS VCCL VCCL sky130_fd_sc_ls__decap_4
XC10 net8 VCCH sky130_fd_pr__cap_mim_m3_1 W=8 L=8 m=1
XC11 net7 VCCH sky130_fd_pr__cap_mim_m3_1 W=16 L=16 m=1
XC12 vbp1 VCCL sky130_fd_pr__cap_mim_m3_1 W=16 L=16 m=1
XC13 vbn1 VSS sky130_fd_pr__cap_mim_m3_1 W=16 L=16 m=1
XC14 VT2 VSS sky130_fd_pr__cap_mim_m3_1 W=16 L=16 m=20
XC15 VT3 VCCL sky130_fd_pr__cap_mim_m3_1 W=16 L=16 m=20
XC16 net12 VCCL sky130_fd_pr__cap_mim_m3_1 W=10 L=10 m=1
XC17 net13 VSS sky130_fd_pr__cap_mim_m3_1 W=10 L=10 m=1
XC18 net14 VCCL sky130_fd_pr__cap_mim_m3_1 W=10 L=10 m=1
XR1 net23 net9 VSS sky130_fd_pr__res_xhigh_po_0p69 L=240 mult=1 m=1
XR7 VSS net23 VSS sky130_fd_pr__res_xhigh_po_0p69 L=240 mult=1 m=1
XM55 net22 net21 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM56 net22 net21 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=2 m=1
XM57 por_h net22 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM58 por_h net22 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=2 m=1
x10 por_h VSS VSS VCCH VCCH porb_h[0] sky130_fd_sc_hvl__inv_16
x8 por_h VSS VSS VCCH VCCH porb_h[1] sky130_fd_sc_hvl__inv_16
Vvgbias net8 ibn180n 0
.save i(vvgbias)
.ends


* expanding   symbol:  EF_LSB_CAP.sym # of pins=9
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_LSB_CAP.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_LSB_CAP.sch
.subckt EF_LSB_CAP VP1 VSS D0 D1 D2 D3 D4 D5 Vref
*.PININFO VP1:B D0:B D1:B D2:B D3:B D4:B VSS:B D5:B Vref:B
XC1 VP1 Vref sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=1
XC2 VP1 D0 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=1
XC6 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=26
XC8 Vref VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=1
XC3 VP1 D1 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=2
XC4 VP1 D2 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=4
XC5 VP1 D3 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=8
XC7 VP1 D4 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=16
XC9 D0 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=1
XC10 D1 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=2
XC11 D2 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=4
XC12 D3 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=8
XC13 D4 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=16
XC14 VSS VSS sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=26
XC15 VP1 D5 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=32
XC16 D5 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=32
.ends


* expanding   symbol:  EF_MSB_CAP.sym # of pins=8
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_MSB_CAP.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_MSB_CAP.sch
.subckt EF_MSB_CAP D8 D10 D9 VP2 D6 VSS D7 D11
*.PININFO D10:B D6:B D7:B D8:B D9:B VP2:B VSS:B D11:B
XC2 D6 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=1
XC3 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=27
XC4 VSS VSS sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=27
XC6 VP2 D6 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=1
XC7 VP2 D7 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=2
XC8 VP2 D8 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=4
XC9 VP2 D9 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=8
XC10 VP2 D10 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=16
XC11 D7 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=2
XC12 D8 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=4
XC13 D9 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=8
XC14 D10 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=16
XC1 VP2 D11 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=32
XC5 D11 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=32
.ends


* expanding   symbol:  EF_SC_CAP.sym # of pins=3
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_SC_CAP.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_SC_CAP.sch
.subckt EF_SC_CAP VP1 VP2 VSS
*.PININFO VP1:B VP2:B VSS:B
XC13 VP1 VP2 sky130_fd_pr__cap_mim_m3_1 W=7 L=7.055 m=1
XC6 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=7 L=7.055 m=9
XC1 VSS VSS sky130_fd_pr__cap_mim_m3_2 W=7 L=7.055 m=9
XC2 VP2 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7.055 m=1
.ends


* expanding   symbol:  EF_AMUX21x.sym # of pins=9
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_AMUX21x.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_AMUX21x.sch
.subckt EF_AMUX21x vdd3p3 vo vss a b sel dvss cm selcm
*.PININFO sel:I vo:B vdd3p3:B vss:B dvss:B a:B b:B cm:B selcm:I
x2 sel dvss dvss vdd3p3 vdd3p3 net1 sky130_fd_sc_hvl__inv_2
x7 selp net2 vss vo a vdd3p3 simple_analog_switch_2
x8 net4 net3 vss vo cm vdd3p3 simple_analog_switch_2
x9 selb net5 vss vo b vdd3p3 simple_analog_switch_2
x11 selp dvss dvss vdd3p3 vdd3p3 net2 sky130_fd_sc_hvl__inv_2
x14 selcm dvss dvss vdd3p3 vdd3p3 net3 sky130_fd_sc_hvl__inv_2
x17 selb dvss dvss vdd3p3 vdd3p3 net5 sky130_fd_sc_hvl__inv_2
x10 net3 dvss dvss vdd3p3 vdd3p3 net4 sky130_fd_sc_hvl__inv_2
x1 selcm net1 dvss dvss vdd3p3 vdd3p3 selb sky130_fd_sc_hvl__nor2_1
x3 sel selcm dvss dvss vdd3p3 vdd3p3 selp sky130_fd_sc_hvl__nor2_1
x4[3] dvss dvss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_8
x4[2] dvss dvss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_8
x4[1] dvss dvss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_8
x4[0] dvss dvss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_8
* noconn dvss
.ends


* expanding   symbol:  simple_analog_switch.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch.sch
.subckt simple_analog_switch on off vss out in vdd
*.PININFO on:I out:B vdd:B vss:B in:B off:I
XM1 in on out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
XM2 in off out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=4 m=1
XM3 out off out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM4 out on out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
XM5 in off in vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM6 in on in vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
.ends


* expanding   symbol:  rheo_column.sym # of pins=13
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rheostat_8bit/xschem/rheo_column.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rheostat_8bit/xschem/rheo_column.sch
.subckt rheo_column b2 b2b b1 b1b b0 b0b vdd dum_in res_in out res_out vss dum_out
*.PININFO res_in:B vss:B vdd:B out:B b0:I b0b:I b1:I b1b:I b2:I b2b:I dum_in:B res_out:B dum_out:B
x1 vdd b0 net8 net1 b0b vss passtrans
x2 vdd b0b net8 net2 b0 vss passtrans
x3 vdd b0 net9 net3 b0b vss passtrans
x4 vdd b0b net9 net4 b0 vss passtrans
x5 vdd b0 net10 net5 b0b vss passtrans
x6 vdd b0b net10 net6 b0 vss passtrans
x7 vdd b0 net11 net7 b0b vss passtrans
x8 vdd b0b net11 res_in b0 vss passtrans
x9 vdd vdd net14 dum_in vss vss passtrans
x10 vdd vdd net15 res_out vss vss passtrans
x11 vdd b1b net13 net11 b1 vss passtrans
x12 vdd b1 net13 net10 b1b vss passtrans
x13 vdd b1b net12 net9 b1 vss passtrans
x14 vdd b1 net12 net8 b1b vss passtrans
x15 vdd b2b out net13 b2 vss passtrans
x16 vdd b2 out net12 b2b vss passtrans
x17 vdd vdd net14 net14 vss vss passtrans
x18 vdd vdd net15 net15 vss vss passtrans
XR1 res_in dum_in sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR2 net7 res_in sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR3 net6 net7 sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR4 net5 net6 sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR5 net4 net5 sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR6 net3 net4 sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR7 net2 net3 sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR8 net1 net2 sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR9 res_out net1 sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
XR10 dum_out res_out sky130_fd_pr__res_generic_po W=0.71 L=2.96 m=1
.ends


* expanding   symbol:  trans_gate.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_vbl_ip__overvoltage/xschem/trans_gate.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_vbl_ip__overvoltage/xschem/trans_gate.sch
.subckt trans_gate in ena_b ena avdd vss out
*.PININFO avdd:B vss:B ena:I ena_b:I in:I out:O
XM1 in ena out vss sky130_fd_pr__nfet_g5v0d10v5 L=5 W=1 nf=1 m=1
XM2 in ena_b out avdd sky130_fd_pr__pfet_g5v0d10v5 L=5 W=6 nf=1 m=1
.ends


* expanding   symbol:  trans_gate_mux.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_vbl_ip__overvoltage/xschem/trans_gate_mux.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_vbl_ip__overvoltage/xschem/trans_gate_mux.sch
.subckt trans_gate_mux in ena_b ena avdd vss out
*.PININFO avdd:B vss:B ena:I ena_b:I in:I out:O
XM1 in ena out vss sky130_fd_pr__nfet_g5v0d10v5 L=3 W=1 nf=1 m=1
XM2 in ena_b out avdd sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1 nf=1 m=1
.ends


* expanding   symbol:  dac_column.sym # of pins=13
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rdac3v_8bit/xschem/dac_column.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__rdac3v_8bit/xschem/dac_column.sch
.subckt dac_column b2 b2b b1 b1b b0 b0b vdd dum_in res_in out res_out vss dum_out
*.PININFO res_in:B vss:B vdd:B out:B b0:I b0b:I b1:I b1b:I b2:I b2b:I dum_in:B res_out:B dum_out:B
x1 vdd b0 net8 net1 b0b vss passtrans
XR1 res_out net1 vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
x2 vdd b0b net8 net2 b0 vss passtrans
x3 vdd b0 net9 net3 b0b vss passtrans
x4 vdd b0b net9 net4 b0 vss passtrans
x5 vdd b0 net10 net5 b0b vss passtrans
x6 vdd b0b net10 net6 b0 vss passtrans
x7 vdd b0 net11 net7 b0b vss passtrans
x8 vdd b0b net11 res_in b0 vss passtrans
x9 vdd vdd net15 dum_in vss vss passtrans
x10 vdd vdd net12 res_out vss vss passtrans
XR2 net1 net2 vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR3 net2 net3 vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR4 net3 net4 vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR5 net4 net5 vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR6 net5 net6 vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR7 net6 net7 vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR9 net7 res_in vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR10 res_in dum_in vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
XR12 dum_out res_out vss sky130_fd_pr__res_high_po_0p35 L=3.16 mult=1 m=1
x11 vdd b1b net14 net11 b1 vss passtrans
x12 vdd b1 net14 net10 b1b vss passtrans
x13 vdd b1b net13 net9 b1 vss passtrans
x14 vdd b1 net13 net8 b1b vss passtrans
x15 vdd b2b out net14 b2 vss passtrans
x16 vdd b2 out net13 b2b vss passtrans
x17 vdd vdd net15 net15 vss vss passtrans
x18 vdd vdd net12 net12 vss vss passtrans
.ends


* expanding   symbol:  isolated_switch_3.sym # of pins=7
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/isolated_switch_3.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/isolated_switch_3.sch
.subckt isolated_switch_3 on off vss out in vdd shunt
*.PININFO on:I out:B vdd:B vss:B in:B off:I shunt:I
XM1 in on net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=12 nf=6 m=1
XM2 in off net1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=24 nf=12 m=1
XM11 net1 on out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=12 nf=6 m=1
XM12 net1 off out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=24 nf=12 m=1
XM17 vss shunt net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends


* expanding   symbol:  isolated_switch_4.sym # of pins=7
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/isolated_switch_4.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__analog_switches/xschem/isolated_switch_4.sch
.subckt isolated_switch_4 on off vss out in vdd shunt
*.PININFO on:I out:B vdd:B vss:B in:B off:I shunt:I
XM1 in on net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=60 nf=6 m=1
XM2 in off net1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=120 nf=12 m=1
XM11 net1 on out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=60 nf=6 m=1
XM12 net1 off out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=120 nf=12 m=1
XM17 vss shunt net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends


* expanding   symbol:  bias_nstack.sym # of pins=5
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/bias_nstack.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/bias_nstack.sch
.subckt bias_nstack itail ena vcasc nbias avss
*.PININFO avss:B ena:I nbias:I itail:B vcasc:B
XM3 net1 nbias avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=1
XM6 vcasc nbias net1 avss sky130_fd_pr__nfet_05v0_nvt L=1 W=3 nf=1 m=1
XM12 itail ena vcasc avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 m=1
XD1 avss ena sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
.ends


* expanding   symbol:  bias_pstack.sym # of pins=7
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/bias_pstack.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/bias_pstack.sch
.subckt bias_pstack avdd pbias pcasc vcasc enb avss itail
*.PININFO avdd:B itail:B enb:I pcasc:I vcasc:B pbias:I avss:B
XM13 net1 pbias avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=3 nf=1 m=1
XM18 itail enb vcasc avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=3 nf=1 m=1
XM14 vcasc pcasc net1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=3 nf=1 m=1
XD1 avss enb sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
.ends


* expanding   symbol:  bias_amp.sym # of pins=7
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/bias_amp.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ef_ip__biasgen/xschem/bias_amp.sch
.subckt bias_amp avdd out inn inp nbias avss ena
*.PININFO inp:I nbias:I inn:I out:O avdd:B avss:B ena:I
XM1 net2 nbias avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM2 out net1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM3 net1 net1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM4 net1 inp vcom avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4 nf=2 m=1
XM5 out inn vcom avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4 nf=2 m=1
XM6 vcom ena net2 avss sky130_fd_pr__nfet_05v0_nvt L=1 W=2 nf=1 m=1
.ends


* expanding   symbol:  rstring_mux.sym # of pins=7
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ajc_ip__brownout/xschem/rstring_mux.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ajc_ip__brownout/xschem/rstring_mux.sch
.subckt rstring_mux avdd vout_brout ena otrip_decoded_avdd[7] otrip_decoded_avdd[6] otrip_decoded_avdd[5] otrip_decoded_avdd[4]
+ otrip_decoded_avdd[3] otrip_decoded_avdd[2] otrip_decoded_avdd[1] otrip_decoded_avdd[0] vtrip_decoded_avdd[7] vtrip_decoded_avdd[6]
+ vtrip_decoded_avdd[5] vtrip_decoded_avdd[4] vtrip_decoded_avdd[3] vtrip_decoded_avdd[2] vtrip_decoded_avdd[1] vtrip_decoded_avdd[0] vout_vunder avss
*.PININFO vout_brout:O otrip_decoded_avdd[7:0]:I vout_vunder:O vtrip_decoded_avdd[7:0]:I ena:I avdd:I avss:I
XR1 net2 net3 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR2 net3 net4 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR0 avss net2 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR3 net4 net5 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR4 net5 net6 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR5 net6 net7 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR6 net7 net8 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR7 net8 net9 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR8 net9 net10 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR9 net10 net11 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR10 net11 net12 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR11 net12 net13 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR12 net13 net14 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR13 net14 net15 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR14 net15 net16 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR15 net16 net17 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR16 net17 net18 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR17 net18 net19 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR18 net19 net20 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR19 net20 net21 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR20 net21 net22 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR21 net22 net23 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR22 net23 net24 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR23 net24 net25 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR24 net25 net26 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR25 net26 net27 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR26 net27 net28 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR27 net28 vtrip7 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR28 vtrip7 vtrip6 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR29 vtrip6 vtrip5 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR30 vtrip5 vtrip4 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR31 vtrip4 vtrip3 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR32 vtrip3 vtrip2 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR33 vtrip2 vtrip1 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR34 vtrip1 vtrip0 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR35 vtrip0 net29 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR36 net29 net30 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR37 net30 net31 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR38 net31 net32 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR39 net32 net33 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR40 net33 net34 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR41 net34 net35 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR42 net35 net36 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR43 net36 net37 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR44 net37 net38 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR45 net38 net39 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR46 net39 net40 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR47 net40 net41 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR48 net41 net42 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR49 net42 net43 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR50 net43 net44 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR51 net44 net45 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR52 net45 net46 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR53 net46 net47 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR54 net47 net48 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR55 net48 net49 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR56 net49 net50 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR57 net50 net51 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR58 net51 net52 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR59 net52 net53 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR60 net53 net54 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR61 net54 net55 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR62 net55 net56 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR63 net56 net57 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR64 net57 net58 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR65 net58 net59 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR66 net59 net60 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR67 net60 net61 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR68 net61 net62 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XR69 net62 net1 avss sky130_fd_pr__res_xhigh_po_1p41 L=35 mult=1 m=1
XMtp[7] vtrip7 otrip_decoded_b_avdd[7] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[6] vtrip6 otrip_decoded_b_avdd[6] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[5] vtrip5 otrip_decoded_b_avdd[5] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[4] vtrip4 otrip_decoded_b_avdd[4] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[3] vtrip3 otrip_decoded_b_avdd[3] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[2] vtrip2 otrip_decoded_b_avdd[2] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[1] vtrip1 otrip_decoded_b_avdd[1] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp[0] vtrip0 otrip_decoded_b_avdd[0] vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[7] vout_brout otrip_decoded_avdd[7] vtrip7 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[6] vout_brout otrip_decoded_avdd[6] vtrip6 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[5] vout_brout otrip_decoded_avdd[5] vtrip5 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[4] vout_brout otrip_decoded_avdd[4] vtrip4 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[3] vout_brout otrip_decoded_avdd[3] vtrip3 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[2] vout_brout otrip_decoded_avdd[2] vtrip2 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[1] vout_brout otrip_decoded_avdd[1] vtrip1 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn[0] vout_brout otrip_decoded_avdd[0] vtrip0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp1[7] vtrip7 vtrip_decoded_b_avdd[7] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp1[6] vtrip6 vtrip_decoded_b_avdd[6] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp1[5] vtrip5 vtrip_decoded_b_avdd[5] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp1[4] vtrip4 vtrip_decoded_b_avdd[4] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp1[3] vtrip3 vtrip_decoded_b_avdd[3] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp1[2] vtrip2 vtrip_decoded_b_avdd[2] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp1[1] vtrip1 vtrip_decoded_b_avdd[1] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtp1[0] vtrip0 vtrip_decoded_b_avdd[0] vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn1[7] vout_vunder vtrip_decoded_avdd[7] vtrip7 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn1[6] vout_vunder vtrip_decoded_avdd[6] vtrip6 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn1[5] vout_vunder vtrip_decoded_avdd[5] vtrip5 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn1[4] vout_vunder vtrip_decoded_avdd[4] vtrip4 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn1[3] vout_vunder vtrip_decoded_avdd[3] vtrip3 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn1[2] vout_vunder vtrip_decoded_avdd[2] vtrip2 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn1[1] vout_vunder vtrip_decoded_avdd[1] vtrip1 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
XMtn1[0] vout_vunder vtrip_decoded_avdd[0] vtrip0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=2
xIinv0[7] otrip_decoded_avdd[7] avss avss avdd avdd otrip_decoded_b_avdd[7] sky130_fd_sc_hvl__inv_1
xIinv0[6] otrip_decoded_avdd[6] avss avss avdd avdd otrip_decoded_b_avdd[6] sky130_fd_sc_hvl__inv_1
xIinv0[5] otrip_decoded_avdd[5] avss avss avdd avdd otrip_decoded_b_avdd[5] sky130_fd_sc_hvl__inv_1
xIinv0[4] otrip_decoded_avdd[4] avss avss avdd avdd otrip_decoded_b_avdd[4] sky130_fd_sc_hvl__inv_1
xIinv0[3] otrip_decoded_avdd[3] avss avss avdd avdd otrip_decoded_b_avdd[3] sky130_fd_sc_hvl__inv_1
xIinv0[2] otrip_decoded_avdd[2] avss avss avdd avdd otrip_decoded_b_avdd[2] sky130_fd_sc_hvl__inv_1
xIinv0[1] otrip_decoded_avdd[1] avss avss avdd avdd otrip_decoded_b_avdd[1] sky130_fd_sc_hvl__inv_1
xIinv0[0] otrip_decoded_avdd[0] avss avss avdd avdd otrip_decoded_b_avdd[0] sky130_fd_sc_hvl__inv_1
xIinv1[7] vtrip_decoded_avdd[7] avss avss avdd avdd vtrip_decoded_b_avdd[7] sky130_fd_sc_hvl__inv_1
xIinv1[6] vtrip_decoded_avdd[6] avss avss avdd avdd vtrip_decoded_b_avdd[6] sky130_fd_sc_hvl__inv_1
xIinv1[5] vtrip_decoded_avdd[5] avss avss avdd avdd vtrip_decoded_b_avdd[5] sky130_fd_sc_hvl__inv_1
xIinv1[4] vtrip_decoded_avdd[4] avss avss avdd avdd vtrip_decoded_b_avdd[4] sky130_fd_sc_hvl__inv_1
xIinv1[3] vtrip_decoded_avdd[3] avss avss avdd avdd vtrip_decoded_b_avdd[3] sky130_fd_sc_hvl__inv_1
xIinv1[2] vtrip_decoded_avdd[2] avss avss avdd avdd vtrip_decoded_b_avdd[2] sky130_fd_sc_hvl__inv_1
xIinv1[1] vtrip_decoded_avdd[1] avss avss avdd avdd vtrip_decoded_b_avdd[1] sky130_fd_sc_hvl__inv_1
xIinv1[0] vtrip_decoded_avdd[0] avss avss avdd avdd vtrip_decoded_b_avdd[0] sky130_fd_sc_hvl__inv_1
xIinv2 ena avss avss avdd avdd ena_b sky130_fd_sc_hvl__inv_1
XMpdn net1 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMpdp avdd ena_b net1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=16
XMdum0 vout_brout avdd vout_brout avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=7
XMdum1 vout_brout avss vout_brout avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=7
XMdum2 vout_brout avdd vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMdum3 vout_vunder avss vout_brout avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMdum4 vout_vunder avdd vout_vunder avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=7
XMdum5 vout_vunder avss vout_vunder avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=7
.ends


* expanding   symbol:  comparator.sym # of pins=7
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ajc_ip__brownout/xschem/comparator.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ajc_ip__brownout/xschem/comparator.sch
.subckt comparator avdd ibias out ena vinn vinp avss
*.PININFO ena:I avdd:I avss:I ibias:I vinn:I vinp:I out:O
XMb vn vn avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMta vt vn avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMl0 vn ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMinv0 ena_b ena avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMinv1 ena_b ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMi0 vnn vinn vt vt sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=16
XMi1 vpp vinp vt vt sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=16
XMld1 vpp vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 m=8
XMh1 vnn vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 m=14
XMh0 vpp vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 m=14
XMld0 vnn vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 m=8
XMpp1 n0 vpp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMnn1 n0 vm avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMpp0 vm vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMnn0 vm vm avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMinv3 n1 n0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 nf=1 m=2
XMinv2 n1 n0 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 nf=1 m=2
XMinv5 out n1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 nf=1 m=8
XMinv4 out n1 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=1 nf=1 m=8
XMl1 vm ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMl3 vnn ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMl4 vpp ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMt1 ibias ena vn avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMt0 vn ena_b ibias avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMl2 n0 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 m=1
XMdum0 vnn avss vt vt sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=16
XMdum1 avss avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1 nf=1 m=4
XMdum2 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 m=2
XMdum3 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=8 W=1 nf=1 m=22
.ends


* expanding   symbol:  ibias_gen.sym # of pins=10
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ajc_ip__brownout/xschem/ibias_gen.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ajc_ip__brownout/xschem/ibias_gen.sch
.subckt ibias_gen avdd ibias0 itest ibias1 ibg_200n vbg_1v2 isrc_sel ena ve avss
*.PININFO vbg_1v2:I ena:I ibias0:O ibg_200n:I isrc_sel:I avdd:I avss:I itest:O ve:I ibias1:O
XM17 vstart vbg_1v2 vn0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=10
XMt9 vstart ena_b vstartena avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMn0 vn0 vn0 ve avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 nf=1 m=2
XMp0 vn0 vp0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 m=2
XMn1 vp0 vn0 vr avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 nf=1 m=2
XMp1 vp0 vp0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 m=2
XMpb0 ibias0 vp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 m=2
XMt0 vp0 isrc_sel vp avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMt1 vp isrc_sel_b vp0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMl6 vp ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMl3 vp0 ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMl1 vn0 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMnn1 vp1 vn1 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=5 nf=1 m=8
XMnn0 vn1 vn1 avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=5 nf=1 m=2
XMl9 vn1 isrc_sel_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMt6 net1 isrc_sel vn1 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMt7 vn1 isrc_sel_b net2 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMpp1 vp1 vp1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 m=2
XMt2 vp isrc_sel_b vp1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMt3 vp1 isrc_sel vp avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMt4 ibg_200n ena net1 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMt5 net2 ena_b ibg_200n avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMl7 vp1 isrc_sel avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMl8 vp1 ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMl10 vn1 ena_b avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMl2 vp0 isrc_sel_b avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMl0 vn0 isrc_sel avss avss sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XMt8 vstartena isrc_sel avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMn2 ena_b ena avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=1
XMp2 ena_b ena avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 m=1
XMn3 isrc_sel_b isrc_sel avss avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=1
XMp3 isrc_sel_b isrc_sel avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 m=1
XMtst itest vp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 m=2
XR1 avss vr avss sky130_fd_pr__res_xhigh_po_1p41 L=700 mult=1 m=1
XMdum0 avss avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=5 nf=1 m=10
XMdum1 vp0 avss vn0 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMdum2 vp avss vp avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMdum3 vp1 avss vn1 avss sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMdum4 ena_b avss isrc_sel_b avss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=1
XMdum5 isrc_sel_b avdd ena_b avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=5 nf=1 m=1
XMdum6 vp0 avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMdum7 vp avdd vp avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMdum8 vn1 avdd vp1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 nf=1 m=1
XMdum9 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 m=4
XMdum10 avss avss ve avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 nf=1 m=1
XMdum11 vr avss ve avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 nf=1 m=1
XMdum12 vr avss avss avss sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 nf=1 m=1
XMpb1 ibias1 vp avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=4 W=5 nf=1 m=2
.ends


* expanding   symbol:  rc_osc.sym # of pins=4
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ajc_ip__brownout/xschem/rc_osc.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ajc_ip__brownout/xschem/rc_osc.sch
.subckt rc_osc dvdd out ena dvss
*.PININFO dvdd:I dvss:I out:O ena:I
XM1 m in dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=2
XM3 m in dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=6
XM2 m n dvss dvss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM4 m n dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=3
XM5 n m dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM6 n m dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=3
XM7 out n dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM8 out n dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=3
XC1 in dvss sky130_fd_pr__cap_mim_m3_2 W=30 L=30 m=6
XR1 net1 in dvss sky130_fd_pr__res_xhigh_po_1p41 L=105 mult=1 m=1
XM12 in ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM9 out ena vr dvss sky130_fd_pr__nfet_01v8 L=0.18 W=1 nf=1 m=1
XM10 out ena_b vr dvdd sky130_fd_pr__pfet_01v8 L=0.18 W=1 nf=1 m=1
XM11 ena_b ena dvss dvss sky130_fd_pr__nfet_01v8 L=0.6 W=1 nf=1 m=1
XM13 ena_b ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.6 W=1 nf=1 m=1
XR2 net2 net1 dvss sky130_fd_pr__res_xhigh_po_1p41 L=105 mult=1 m=1
XR3 net3 net2 dvss sky130_fd_pr__res_xhigh_po_1p41 L=105 mult=1 m=1
XR4 net4 net3 dvss sky130_fd_pr__res_xhigh_po_1p41 L=105 mult=1 m=1
XR5 net5 net4 dvss sky130_fd_pr__res_xhigh_po_1p41 L=105 mult=1 m=1
XR6 net6 net5 dvss sky130_fd_pr__res_xhigh_po_1p41 L=105 mult=1 m=1
XR7 net7 net6 dvss sky130_fd_pr__res_xhigh_po_1p41 L=105 mult=1 m=1
XR8 net8 net7 dvss sky130_fd_pr__res_xhigh_po_1p41 L=105 mult=1 m=1
XR9 net9 net8 dvss sky130_fd_pr__res_xhigh_po_1p41 L=105 mult=1 m=1
XR10 vr net9 dvss sky130_fd_pr__res_xhigh_po_1p41 L=105 mult=1 m=1
XMdum0 vr dvss dvss dvss sky130_fd_pr__nfet_01v8 L=0.6 W=1 nf=1 m=1
XMdum1 out dvss dvss dvss sky130_fd_pr__nfet_01v8 L=0.18 W=1 nf=1 m=1
XMdum2 m dvss dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XMdum3 n dvss dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XMdum4 m dvdd n dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=1
XMdum5 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.18 W=1 nf=1 m=1
XMdum6 ena_b dvdd vr dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=1
XMdum7 dvdd dvdd out dvdd sky130_fd_pr__pfet_01v8 L=0.18 W=1 nf=1 m=1
.ends


* expanding   symbol:  schmitt_trigger.sym # of pins=4
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_ajc_ip__brownout/xschem/schmitt_trigger.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_ajc_ip__brownout/xschem/schmitt_trigger.sch
.subckt schmitt_trigger dvdd in out dvss
*.PININFO dvdd:I dvss:I out:O in:I
XM1 m in dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=2
XM3 m in dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=6
XM2 m out dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM4 m out dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=3
XM5 out m dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XM6 out m dvdd dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=3
XMdum0 m dvss dvss dvss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 m=1
XMdum1 dvdd dvdd m dvdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 m=1
.ends


* expanding   symbol:  Universal_R_2R_Block2.sym # of pins=9
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/Universal_R_2R_Block2.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/Universal_R_2R_Block2.sch
.subckt Universal_R_2R_Block2 VD DVDD VIRTOUT CMOUT R2RIN R2ROUT DVSS AVDD AVSS
*.PININFO VD:B R2ROUT:B R2RIN:B VIRTOUT:B CMOUT:B DVDD:B AVSS:B AVDD:B DVSS:B
.save v(vx)
x12 net6 VDBAR VDbuf VX AVSS AVDD T_Gate_5V
x13 net5 VDbuf VDBAR VX AVSS AVDD T_Gate_5V
VI12 net1 net4 0
.save i(vi12)
VI1 net1 R2ROUT 0
.save i(vi1)
.save v(vdbar)
.save v(vdbuf)
VI2 net5 CMOUT 0
.save i(vi2)
VI3 net6 VIRTOUT 0
.save i(vi3)
VI4 R2RIN net2 0
.save i(vi4)
x1 VD DVDD DVSS DVSS AVDD AVDD VDbuf sky130_fd_sc_hvl__lsbuflv2hv_1
x2 VDbuf DVSS DVSS AVDD AVDD VDBAR sky130_fd_sc_hvl__inv_1
XR1 net4 net3 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=20 mult=1 m=1
XR3 net3 VX AVSS sky130_fd_pr__res_xhigh_po_0p35 L=20 mult=1 m=1
XR2 net1 net2 AVSS sky130_fd_pr__res_xhigh_po_0p35 L=20 mult=1 m=1
x3 VD DVSS DVSS AVDD AVDD sky130_fd_sc_hvl__diode_2
.ends


* expanding   symbol:  Output_OA.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/Output_OA.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/Output_OA.sch
.subckt Output_OA VDD VOUT VINN VINP VBIAS VSS
*.PININFO VINN:B VINP:B VOUT:B VDD:B VSS:B VBIAS:B
XM1 net4 VINN net1 net1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7.5 nf=1 m=1
XM2 net3 VINP net1 net1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7.5 nf=1 m=1
VISink net1 net2 0
.save i(visink)
XM6 net5 net5 net6 net6 sky130_fd_pr__pfet_01v8_lvt L=5 W=20 nf=1 m=2
XM7 net7 net5 net6 net6 sky130_fd_pr__pfet_01v8_lvt L=5 W=20 nf=1 m=2
VD1 net5 net8 0
.save i(vd1)
VID2 net7 net9 0
.save i(vid2)
VID1 VOUT net12 0
.save i(vid1)
VID3 net11 VOUT 0
.save i(vid3)
.save v(vinn)
.save v(vinp)
.save v(vout)
VIBIAS VBIAS net10 0
.save i(vibias)
XM10 net8 VINN net4 net4 sky130_fd_pr__nfet_05v0_nvt L=2 W=1 nf=1 m=25
XM12 net9 VINP net3 net3 sky130_fd_pr__nfet_05v0_nvt L=2 W=1 nf=1 m=25
XM3 net2 net10 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=20
XM5 net12 net10 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=200
XM8 net11 net7 net6 net6 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 m=10
VIVDD VDD net6 0
.save i(vivdd)
XC1 net7 net13 sky130_fd_pr__cap_mim_m3_1 W=10 L=10 m=15
XR1 net13 VOUT VSS sky130_fd_pr__res_high_po_0p69 L=41 mult=1 m=1
.ends


* expanding   symbol:  x1_x32_OA.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/x1_x32_OA.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/x1_x32_OA.sch
.subckt x1_x32_OA VDD VOUT VINN VINP VBIAS VSS
*.PININFO VINN:B VINP:B VOUT:B VDD:B VSS:B VBIAS:B
XM1 net4 VINN net1 net1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7.5 nf=1 m=1
XM2 net3 VINP net1 net1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7.5 nf=1 m=1
VISink net1 net2 0
.save i(visink)
XM6 net5 net5 net6 net6 sky130_fd_pr__pfet_01v8_lvt L=5 W=20 nf=1 m=2
XM7 net7 net5 net6 net6 sky130_fd_pr__pfet_01v8_lvt L=5 W=20 nf=1 m=2
VD1 net5 net8 0
.save i(vd1)
VID2 net7 net9 0
.save i(vid2)
VID1 VOUT net12 0
.save i(vid1)
VID3 net11 VOUT 0
.save i(vid3)
.save v(vinn)
.save v(vinp)
.save v(vout)
VIBIAS VBIAS net10 0
.save i(vibias)
XM10 net8 VINN net4 net4 sky130_fd_pr__nfet_05v0_nvt L=2 W=1 nf=1 m=25
XM12 net9 VINP net3 net3 sky130_fd_pr__nfet_05v0_nvt L=2 W=1 nf=1 m=25
XM3 net2 net10 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=15
XM5 net12 net10 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=100
XM8 net11 net7 net6 net6 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 m=10
VIVDD VDD net6 0
.save i(vivdd)
XC1 net7 net13 sky130_fd_pr__cap_mim_m3_1 W=10 L=10 m=15
XR1 net13 VOUT VSS sky130_fd_pr__res_high_po_0p69 L=41 mult=1 m=1
.ends


* expanding   symbol:  Input_Stage_OA1.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/Input_Stage_OA1.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/Input_Stage_OA1.sch
.subckt Input_Stage_OA1 VDD VOUT VINN VINP VBIAS VSS
*.PININFO VINN:B VINP:B VOUT:B VDD:B VSS:B VBIAS:B
XM1 net4 VINN net1 net1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7.5 nf=1 m=1
XM2 net3 VINP net1 net1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7.5 nf=1 m=1
VISink net1 net2 0
.save i(visink)
XM6 net5 net5 net6 net6 sky130_fd_pr__pfet_01v8_lvt L=5 W=20 nf=1 m=2
XM7 net7 net5 net6 net6 sky130_fd_pr__pfet_01v8_lvt L=5 W=20 nf=1 m=2
VD1 net5 net8 0
.save i(vd1)
VID2 net7 net9 0
.save i(vid2)
VID1 VOUT net12 0
.save i(vid1)
VID3 net11 VOUT 0
.save i(vid3)
.save v(vinn)
.save v(vinp)
.save v(vout)
VIBIAS VBIAS net10 0
.save i(vibias)
XM10 net8 VINN net4 net4 sky130_fd_pr__nfet_05v0_nvt L=2 W=1 nf=1 m=25
XM12 net9 VINP net3 net3 sky130_fd_pr__nfet_05v0_nvt L=2 W=1 nf=1 m=25
XM3 net2 net10 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=10
XM5 net12 net10 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=20
XM8 net11 net7 net6 net6 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 m=10
VIVDD VDD net6 0
.save i(vivdd)
XC1 net7 net13 sky130_fd_pr__cap_mim_m3_1 W=10 L=10 m=15
XR2 net13 VOUT VSS sky130_fd_pr__res_high_po_0p69 L=41 mult=1 m=1
.ends


* expanding   symbol:  Input_Stage_OA2.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/Input_Stage_OA2.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/Input_Stage_OA2.sch
.subckt Input_Stage_OA2 VDD VOUT VINN VINP VBIAS VSS
*.PININFO VINN:B VINP:B VOUT:B VDD:B VSS:B VBIAS:B
XM1 net4 VINN net1 net1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7.5 nf=1 m=1
XM2 net3 VINP net1 net1 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=7.5 nf=1 m=1
VISink net1 net2 0
.save i(visink)
XM6 net5 net5 net6 net6 sky130_fd_pr__pfet_01v8_lvt L=5 W=20 nf=1 m=2
XM7 net7 net5 net6 net6 sky130_fd_pr__pfet_01v8_lvt L=5 W=20 nf=1 m=2
VD1 net5 net8 0
.save i(vd1)
VID2 net7 net9 0
.save i(vid2)
VID1 VOUT net12 0
.save i(vid1)
VID3 net11 VOUT 0
.save i(vid3)
.save v(vinn)
.save v(vinp)
.save v(vout)
VIBIAS VBIAS net10 0
.save i(vibias)
XM10 net8 VINN net4 net4 sky130_fd_pr__nfet_05v0_nvt L=2 W=1 nf=1 m=25
XM12 net9 VINP net3 net3 sky130_fd_pr__nfet_05v0_nvt L=2 W=1 nf=1 m=25
XM3 net2 net10 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=20
XM5 net12 net10 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=5 nf=1 m=100
XM8 net11 net7 net6 net6 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 m=10
VIVDD VDD net6 0
.save i(vivdd)
XC1 net7 net13 sky130_fd_pr__cap_mim_m3_1 W=10 L=10 m=15
XR1 net13 VOUT VSS sky130_fd_pr__res_high_po_0p69 L=41 mult=1 m=1
.ends


* expanding   symbol:  bandgap/bg_res.sym # of pins=5
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_cw_ip/xschem/bandgap/bg_res.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_cw_ip/xschem/bandgap/bg_res.sch
.subckt bg_res b a d c vss
*.PININFO a:I b:I c:O d:O vss:B
XR1 net1 a vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR2 net2 b vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR3 net6 net1 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR4 net5 net2 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR5 net3 net6 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR6 net4 net5 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR7 net10 net3 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR8 net9 net4 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR9 net7 net10 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR10 net8 net9 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR11 net12 net7 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR12 net11 net8 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR13 net14 net12 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR14 net13 net11 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR15 net16 net14 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR16 net15 net13 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR17 net18 net16 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR18 net17 net15 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR19 c net18 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
XR20 d net17 vss sky130_fd_pr__res_xhigh_po_0p69 L=13 mult=1 m=1
.ends


* expanding   symbol:  bandgap/bg_trim.sym # of pins=4
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_cw_ip/xschem/bandgap/bg_trim.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_cw_ip/xschem/bandgap/bg_trim.sch
.subckt bg_trim top bot ctl[15] ctl[14] ctl[13] ctl[12] ctl[11] ctl[10] ctl[9] ctl[8] ctl[7] ctl[6] ctl[5] ctl[4] ctl[3] ctl[2]
+ ctl[1] ctl[0] vss
*.PININFO vss:B ctl[15:0]:I bot:B top:B
XM0 net1 ctl[0] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM1 net2 ctl[1] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM2 net3 ctl[2] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM3 net4 ctl[3] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM4 net5 ctl[4] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM5 net6 ctl[5] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM6 net7 ctl[6] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM7 net8 ctl[7] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM12 net10 ctl[12] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM13 net11 ctl[13] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM14 net12 ctl[14] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM15 top ctl[15] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM8 net13 ctl[8] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM9 net14 ctl[9] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM10 net15 ctl[10] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XM11 net9 ctl[11] bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 m=1
XR15 net12 top vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR1 net1 net2 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR16 bot net1 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR2 net2 net3 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR3 net3 net4 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR4 net4 net5 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR5 net5 net6 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR6 net6 net7 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR7 net7 net8 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR8 net8 net13 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR9 net13 net14 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR10 net14 net15 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR11 net15 net9 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR12 net9 net10 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR13 net10 net11 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
XR14 net11 net12 vss sky130_fd_pr__res_high_po_1p41 L=2.92 mult=1 m=1
.ends


* expanding   symbol:  opamp/se_folded_cascode_p.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_cw_ip/xschem/opamp/se_folded_cascode_p.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_cw_ip/xschem/opamp/se_folded_cascode_p.sch
.subckt se_folded_cascode_p vdd out inp inn vss bias
*.PININFO inn:I inp:I out:O bias:B vdd:B vss:B
XM3 out1p inn diff vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 m=8
XM2 out1n inp diff vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 m=8
XM1 diff vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=16
XM4 out1n vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=16
XM5 out1p vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=16
XM6 mirr vbn2 out1n vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=8
XM7 out vbn2 out1p vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=8
XM8 mirr bias nd10 vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=8
XM9 out bias nd11 vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=8
XM10 nd10 mirr vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=8
XM11 nd11 mirr vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=8
XMB1 bias bias vbp1 vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=4
XMB2 vbp1 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=4
XMB3 vbn2 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=4
XMB4 vbn2 vbn2 vbn1 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=4
XMB5 vbn1 vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=4
XMDUM1[43] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[42] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[41] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[40] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[39] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[38] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[37] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[36] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[35] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[34] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[33] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[32] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[31] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[30] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[29] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[28] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[27] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[26] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[25] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[24] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[23] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[22] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[21] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[20] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[19] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[18] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[17] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[16] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[15] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[14] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[13] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[12] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[11] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[10] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[9] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[8] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[7] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[6] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[5] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[4] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[3] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[2] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[1] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM1[0] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM2[3] mirr mirr mirr vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM2[2] mirr mirr mirr vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM2[1] mirr mirr mirr vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM2[0] mirr mirr mirr vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM3[3] bias bias bias vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM3[2] bias bias bias vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM3[1] bias bias bias vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM3[0] bias bias bias vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 m=1
XMDUM4[23] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[22] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[21] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[20] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[19] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[18] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[17] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[16] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[15] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[14] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[13] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[12] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[11] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[10] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[9] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[8] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[7] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[6] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[5] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[4] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[3] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[2] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[1] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM4[0] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM5[3] vbn2 vbn2 vbn2 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM5[2] vbn2 vbn2 vbn2 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM5[1] vbn2 vbn2 vbn2 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM5[0] vbn2 vbn2 vbn2 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 m=1
XMDUM6[43] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[42] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[41] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[40] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[39] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[38] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[37] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[36] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[35] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[34] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[33] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[32] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[31] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[30] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[29] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[28] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[27] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[26] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[25] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[24] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[23] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[22] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[21] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[20] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[19] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[18] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[17] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[16] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[15] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[14] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[13] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[12] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[11] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[10] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[9] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[8] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[7] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[6] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[5] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[4] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[3] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[2] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[1] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM6[0] vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM7[3] diff diff diff vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 m=1
XMDUM7[2] diff diff diff vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 m=1
XMDUM7[1] diff diff diff vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 m=1
XMDUM7[0] diff diff diff vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 m=1
XMDUM8[31] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[30] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[29] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[28] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[27] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[26] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[25] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[24] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[23] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[22] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[21] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[20] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[19] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[18] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[17] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[16] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[15] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[14] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[13] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[12] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[11] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[10] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[9] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[8] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[7] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[6] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[5] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[4] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[3] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[2] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[1] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XMDUM8[0] vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
.ends


* expanding   symbol:  levelShifter.sym # of pins=5
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_sw_ip__por/xschem/levelShifter.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_sw_ip__por/xschem/levelShifter.sch
.subckt levelShifter ain aout VCCL VSS VCCH
*.PININFO VCCL:I VSS:I ain:I aout:O VCCH:I
XM12 net1 S1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3.6 nf=1 m=1
XM13 aob net1 VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5.8 nf=2 m=1
XM6 S1 ain VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM1 S1 ain VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
XM2 net1 aob VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5.8 nf=2 m=1
XM3 aob S1B VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3.6 nf=1 m=1
XM4 S1B S1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM5 S1B S1 VCCL VCCL sky130_fd_pr__pfet_01v8 L=0.15 W=1.4 nf=2 m=1
XM7 aout aob VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1.8 nf=1 m=1
XM8 aout aob VCCH VCCH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5.8 nf=2 m=1
XC1 VCCH aob sky130_fd_pr__cap_mim_m3_1 W=2 L=2 m=1
.ends


* expanding   symbol:  TieH_1p8.sym # of pins=3
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_sw_ip__por/xschem/TieH_1p8.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_sw_ip__por/xschem/TieH_1p8.sch
.subckt TieH_1p8 TieH VSS VCC
*.PININFO VCC:I VSS:I TieH:B
XM4 net1 net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 m=1
XM5 TieH net1 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=2 m=1
.ends


* expanding   symbol:  T_Gate_5V.sym # of pins=6
** sym_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/T_Gate_5V.sym
** sch_path: /home/tim/gits/frigate_analog/dependencies/sky130_pa_ip__instramp/xschem/T_Gate_5V.sch
.subckt T_Gate_5V UPPER PGATE NGATE LOWER AVSS AVDD
*.PININFO PGATE:B UPPER:B LOWER:B NGATE:B AVDD:B AVSS:B
VI6 net2 net1 0
.save i(vi6)
VI1 net2 net3 0
.save i(vi1)
VI2 net6 net4 0
.save i(vi2)
VI3 net5 net4 0
.save i(vi3)
XM1 net5 net7 net1 AVSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM2 net3 net8 net6 AVDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
VI4 net4 UPPER 0
.save i(vi4)
VI5 LOWER net2 0
.save i(vi5)
VI7 PGATE net8 0
.save i(vi7)
VI8 net7 NGATE 0
.save i(vi8)
.ends

.end
