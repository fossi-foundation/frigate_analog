magic
tech sky130A
magscale 1 2
timestamp 1723666764
<< psubdiff >>
rect 30081 20698 30105 21096
rect 40871 20698 40895 21096
<< psubdiffcont >>
rect 30105 20698 40871 21096
<< locali >>
rect 30054 21096 40924 21132
rect 30054 20698 30105 21096
rect 40871 20698 40924 21096
rect 30054 20674 40924 20698
<< viali >>
rect 30105 20698 40871 21096
<< metal1 >>
rect 36393 25005 47925 25017
rect 36393 24953 36420 25005
rect 36592 24953 47925 25005
rect 36393 24947 47925 24953
rect 3566 24059 33342 24073
rect 3566 24007 33164 24059
rect 33336 24007 33342 24059
rect 3566 23986 33342 24007
rect 3566 23449 3653 23986
rect 4278 23850 33790 23866
rect 4278 23798 33612 23850
rect 33784 23798 33790 23850
rect 4278 23779 33790 23798
rect 4278 23384 4365 23779
rect 23920 23630 36030 23646
rect 23920 23578 35852 23630
rect 36024 23578 36030 23630
rect 23920 23563 36030 23578
rect 23920 23419 24003 23563
rect 29701 23208 30104 23221
rect 29701 22941 29714 23208
rect 29692 22830 29714 22941
rect 30092 22830 30104 23208
rect 29692 22818 30104 22830
rect 40768 23089 41174 23101
rect 29692 22141 30092 22818
rect 40768 22711 40783 23089
rect 41161 22711 41174 23089
rect 40768 22696 41174 22711
rect 29418 21965 30092 22141
rect 25596 21390 26513 21401
rect 25596 21160 25614 21390
rect 25782 21160 26513 21390
rect 25596 21151 26513 21160
rect 29714 21138 30092 21965
rect 40783 21138 41161 22696
rect 82548 21505 83376 22331
rect 26252 21066 26639 21123
rect 29714 21096 41161 21138
rect 26252 18647 26309 21066
rect 29714 20698 30105 21096
rect 40871 20698 41161 21096
rect 29714 20629 41161 20698
rect 29714 20587 30092 20629
rect 29261 20337 30092 20587
rect 26532 18796 26962 18856
rect 26532 18647 26592 18796
rect 26252 18590 26592 18647
rect 26532 18488 26592 18590
rect 26894 18488 26962 18796
rect 26532 18426 26962 18488
rect 27262 18310 27530 19708
rect 25600 18296 27530 18310
rect 25600 18060 25614 18296
rect 25780 18060 27530 18296
rect 25600 18042 27530 18060
rect 29714 13282 30092 20337
rect 31769 18580 32287 18595
rect 31769 18091 31784 18580
rect 32273 18091 32287 18580
rect 31769 18074 32287 18091
rect 31784 13171 32273 18074
rect 40783 14562 41161 20629
rect 43156 18862 43569 18875
rect 43156 18484 43174 18862
rect 43552 18484 43569 18862
rect 43156 18469 43569 18484
rect 43174 14562 43552 18469
<< via1 >>
rect 36420 24953 36592 25005
rect 33164 24007 33336 24059
rect 33612 23798 33784 23850
rect 35852 23578 36024 23630
rect 29714 22830 30092 23208
rect 40783 22711 41161 23089
rect 25614 21160 25782 21390
rect 26592 18488 26894 18796
rect 25614 18060 25780 18296
rect 31784 18091 32273 18580
rect 43174 18484 43552 18862
<< metal2 >>
rect 1966 24066 2385 24071
rect 1966 23666 1976 24066
rect 2376 23666 2385 24066
rect 1966 23662 2385 23666
rect 819 23452 1884 23467
rect 1976 23461 2376 23662
rect 6366 23519 6375 23919
rect 6775 23519 8274 23919
rect 7874 23461 8274 23519
rect 9774 23790 10174 23813
rect 819 23081 838 23452
rect 1303 23081 1884 23452
rect 9774 23427 9792 23790
rect 10155 23427 10174 23790
rect 11121 23567 26188 23714
rect 11121 23440 11268 23567
rect 9774 23409 10174 23427
rect 819 23066 1884 23081
rect 25600 21390 25798 21412
rect 25600 21160 25614 21390
rect 25782 21160 25798 21390
rect 25600 18296 25798 21160
rect 25600 18060 25614 18296
rect 25780 18060 25798 18296
rect 25600 5452 25798 18060
rect 25502 5390 25884 5452
rect 25502 4474 25564 5390
rect 25826 4474 25884 5390
rect 25502 4406 25884 4474
rect 26041 1692 26188 23567
rect 29701 23208 30104 23221
rect 29701 22830 29714 23208
rect 30092 22830 30104 23208
rect 29701 22818 30104 22830
rect 31504 22582 31532 25600
rect 26600 22554 31532 22582
rect 31952 19446 31980 25600
rect 29298 19418 31980 19446
rect 26532 18796 26962 18856
rect 26532 18488 26592 18796
rect 26894 18488 26962 18796
rect 26532 18426 26962 18488
rect 31769 18580 32287 18595
rect 31769 18091 31784 18580
rect 32273 18091 32287 18580
rect 31769 18074 32287 18091
rect 32400 14210 32428 25600
rect 32848 15085 32876 25600
rect 33296 24065 33324 25600
rect 33164 24059 33336 24065
rect 33164 24001 33336 24007
rect 33744 23856 33772 25600
rect 34192 24069 34220 25600
rect 34176 24060 34356 24069
rect 34176 23991 34356 24000
rect 34640 23945 34668 25600
rect 34624 23936 34804 23945
rect 34624 23867 34804 23876
rect 33612 23850 33784 23856
rect 33612 23792 33784 23798
rect 32832 15076 32992 15085
rect 32832 15007 32992 15016
rect 31333 14182 32428 14210
rect 30504 14064 30668 14073
rect 30504 14008 30512 14064
rect 30504 13999 30668 14008
rect 30504 13736 30549 13999
rect 31333 13733 31378 14182
rect 35088 14075 35116 25600
rect 35536 15395 35564 25600
rect 35984 23636 36012 25600
rect 36432 25011 36460 25600
rect 36420 25005 36592 25011
rect 36420 24947 36592 24953
rect 35852 23630 36024 23636
rect 35852 23572 36024 23578
rect 40768 23089 41174 23101
rect 40768 22711 40783 23089
rect 41161 22711 41174 23089
rect 40768 22696 41174 22711
rect 82548 21505 83376 22331
rect 43156 18862 43569 18875
rect 43156 18484 43174 18862
rect 43552 18484 43569 18862
rect 43156 18469 43569 18484
rect 35536 15367 41820 15395
rect 41775 14919 41820 15367
rect 42504 15074 42681 15083
rect 42680 15018 42681 15074
rect 42504 15009 42681 15018
rect 42636 14919 42681 15009
rect 34932 14066 35132 14075
rect 34932 13997 35132 14006
rect 33458 9667 34404 9722
rect 33458 8013 33545 9667
rect 34317 8013 34404 9667
rect 33458 7910 34404 8013
rect 44943 9627 46398 9715
rect 44943 8021 45015 9627
rect 46295 8021 46398 9627
rect 44943 7925 46398 8021
rect 27733 5627 28735 5699
rect 27733 4029 27804 5627
rect 28679 4029 28735 5627
rect 27733 3950 28735 4029
rect 38097 5627 39751 5699
rect 38097 4021 38176 5627
rect 39679 4021 39751 5627
rect 38097 3942 39751 4021
rect 26041 1679 26388 1692
rect 26041 1523 26388 1532
rect 20506 400 20710 620
rect 9000 196 20710 400
rect 22966 400 23170 688
rect 68513 516 69015 628
rect 22966 196 31300 400
rect 9000 0 9300 196
rect 31000 0 31300 196
rect 53000 300 69015 516
rect 69512 300 69513 628
rect 69525 311 69993 612
rect 70015 300 75300 516
rect 53000 0 53300 300
rect 75000 0 75300 300
<< via2 >>
rect 1976 23666 2376 24066
rect 6375 23519 6775 23919
rect 838 23081 1303 23452
rect 9792 23427 10155 23790
rect 25564 4474 25826 5390
rect 29714 22830 30092 23208
rect 26592 18488 26894 18796
rect 31784 18091 32273 18580
rect 34176 24000 34356 24060
rect 34624 23876 34804 23936
rect 32832 15016 32992 15076
rect 30512 14008 30668 14064
rect 40783 22711 41161 23089
rect 43174 18484 43552 18862
rect 42504 15018 42680 15074
rect 34932 14006 35132 14066
rect 33545 8013 34317 9667
rect 45015 8021 46295 9627
rect 27804 4029 28679 5627
rect 38176 4021 39679 5627
rect 26041 1532 26388 1679
<< metal3 >>
rect 50993 25423 82195 25483
rect 1971 24066 2381 24071
rect 95 23666 101 24066
rect 591 23666 1976 24066
rect 2376 23666 2381 24066
rect 34171 24062 34361 24065
rect 50993 24062 51053 25423
rect 34171 24060 51053 24062
rect 34171 24000 34176 24060
rect 34356 24002 51053 24060
rect 51113 25269 80875 25329
rect 82135 25318 82195 25423
rect 34356 24000 34361 24002
rect 34171 23995 34361 24000
rect 51113 23941 51173 25269
rect 34619 23936 51173 23941
rect 1971 23661 2381 23666
rect 6361 23924 6788 23930
rect 6361 23514 6370 23924
rect 6780 23514 6788 23924
rect 34619 23876 34624 23936
rect 34804 23881 51173 23936
rect 34804 23876 34809 23881
rect 34619 23871 34809 23876
rect 6361 23507 6788 23514
rect 9774 23790 10174 23809
rect 819 23452 1321 23467
rect 819 23081 838 23452
rect 1303 23081 1321 23452
rect 9774 23427 9792 23790
rect 10155 23427 10174 23790
rect 9774 23409 10174 23427
rect 82558 23579 83392 23617
rect 819 23066 1321 23081
rect 29701 23213 30104 23221
rect 29701 22825 29709 23213
rect 30097 22825 30104 23213
rect 29701 22818 30104 22825
rect 40768 23094 41174 23101
rect 40768 22706 40778 23094
rect 41166 22706 41174 23094
rect 82558 22795 82573 23579
rect 83368 22795 83392 23579
rect 82558 22766 83392 22795
rect 40768 22696 41174 22706
rect 82548 22319 83376 22331
rect 82548 21519 82565 22319
rect 83365 21519 83376 22319
rect 82548 21505 83376 21519
rect 82565 19233 83365 20928
rect 43156 18867 43569 18875
rect 26532 18796 26962 18856
rect 26532 18488 26592 18796
rect 26894 18488 26962 18796
rect 26532 18426 26962 18488
rect 31769 18585 32287 18595
rect 31769 18086 31779 18585
rect 32278 18086 32287 18585
rect 43156 18479 43169 18867
rect 43557 18479 43569 18867
rect 43156 18469 43569 18479
rect 82565 18427 83365 18433
rect 31769 18074 32287 18086
rect 32827 15076 32997 15081
rect 42499 15076 42685 15079
rect 32827 15016 32832 15076
rect 32992 15074 42685 15076
rect 32992 15018 42504 15074
rect 42680 15018 42685 15074
rect 32992 15016 42685 15018
rect 32827 15011 32997 15016
rect 42499 15013 42685 15016
rect 30507 14066 30673 14069
rect 34927 14066 35137 14071
rect 30507 14064 34932 14066
rect 30507 14008 30512 14064
rect 30668 14008 34932 14064
rect 30507 14006 34932 14008
rect 35132 14006 35137 14066
rect 30507 14003 30673 14006
rect 34927 14001 35137 14006
rect 33458 9667 34404 9722
rect 33458 8013 33545 9667
rect 34317 8013 34404 9667
rect 33458 7910 34404 8013
rect 44943 9627 46398 9715
rect 44943 8021 45015 9627
rect 46295 8021 46398 9627
rect 82565 9357 83365 10029
rect 82565 8551 83365 8557
rect 44943 7925 46398 8021
rect 27733 5627 28735 5699
rect 25502 5390 25884 5452
rect 25502 4474 25564 5390
rect 25826 4474 25884 5390
rect 25502 4406 25884 4474
rect 27733 4029 27804 5627
rect 28679 4029 28735 5627
rect 27733 3950 28735 4029
rect 38097 5627 39751 5699
rect 38097 4021 38176 5627
rect 39679 4021 39751 5627
rect 38097 3942 39751 4021
rect 82565 5045 83365 5051
rect 82565 3527 83365 4245
rect 26036 1679 26393 1684
rect 26036 1532 26041 1679
rect 26388 1532 46491 1679
rect 26036 1527 26393 1532
rect 46344 959 46491 1532
rect 46344 954 46697 959
rect 46691 807 46697 954
rect 78024 824 78652 1003
rect 79231 824 79237 1003
rect 46344 801 46697 807
<< via3 >>
rect 101 23666 591 24066
rect 6370 23919 6780 23924
rect 6370 23519 6375 23919
rect 6375 23519 6775 23919
rect 6775 23519 6780 23919
rect 6370 23514 6780 23519
rect 838 23081 1303 23452
rect 9792 23427 10155 23790
rect 29709 23208 30097 23213
rect 29709 22830 29714 23208
rect 29714 22830 30092 23208
rect 30092 22830 30097 23208
rect 29709 22825 30097 22830
rect 40778 23089 41166 23094
rect 40778 22711 40783 23089
rect 40783 22711 41161 23089
rect 41161 22711 41166 23089
rect 40778 22706 41166 22711
rect 82573 22795 83368 23579
rect 82565 21519 83365 22319
rect 26592 18488 26894 18796
rect 31779 18580 32278 18585
rect 31779 18091 31784 18580
rect 31784 18091 32273 18580
rect 32273 18091 32278 18580
rect 31779 18086 32278 18091
rect 43169 18862 43557 18867
rect 43169 18484 43174 18862
rect 43174 18484 43552 18862
rect 43552 18484 43557 18862
rect 43169 18479 43557 18484
rect 82565 18433 83365 19233
rect 33545 8013 34317 9667
rect 45015 8021 46295 9627
rect 82565 8557 83365 9357
rect 25564 4474 25826 5390
rect 27804 4029 28679 5627
rect 38176 4021 39679 5627
rect 82565 4245 83365 5045
rect 46344 807 46691 954
rect 78652 824 79231 1003
<< metal4 >>
rect 98 24066 598 24077
rect 98 23666 101 24066
rect 591 23666 598 24066
rect 98 5814 598 23666
rect 6369 23924 6781 23925
rect 6369 23514 6370 23924
rect 6780 23514 6781 23924
rect 6369 23513 6781 23514
rect 9774 23790 10174 23809
rect 819 23452 1321 23467
rect 819 23081 838 23452
rect 1303 23081 1321 23452
rect 819 23066 1321 23081
rect 820 9780 1320 23066
rect 6375 19797 6614 23513
rect 9774 23427 9792 23790
rect 10155 23427 10174 23790
rect 9774 23409 10174 23427
rect 82558 23579 83392 23617
rect 26778 23264 27188 23288
rect 26778 22916 26800 23264
rect 27164 22916 27188 23264
rect 26778 22890 27188 22916
rect 29701 23214 30104 23221
rect 26778 21680 26958 22890
rect 29701 22824 29708 23214
rect 30098 22824 30104 23214
rect 29701 22818 30104 22824
rect 40768 23095 41174 23101
rect 40768 22705 40777 23095
rect 41167 22705 41174 23095
rect 82558 22795 82573 23579
rect 83368 22795 83392 23579
rect 82558 22766 83392 22795
rect 40768 22696 41174 22705
rect 82548 22320 83376 22331
rect 82548 21518 82564 22320
rect 83366 21518 83376 22320
rect 82548 21505 83376 21518
rect 6375 19773 6919 19797
rect 6375 17856 6405 19773
rect 6891 17856 6919 19773
rect 43156 18868 43569 18875
rect 26532 18796 26962 18856
rect 26532 18488 26592 18796
rect 26894 18488 26962 18796
rect 26532 18426 26962 18488
rect 31769 18586 32287 18595
rect 31769 18085 31778 18586
rect 32279 18085 32287 18586
rect 43156 18478 43168 18868
rect 43558 18478 43569 18868
rect 43156 18469 43569 18478
rect 31769 18074 32287 18085
rect 6375 17826 6919 17856
rect 820 7841 846 9780
rect 1276 7841 1320 9780
rect 820 7809 1320 7841
rect 25670 17396 26216 17478
rect 25670 16042 25734 17396
rect 26134 16042 26216 17396
rect 25670 9724 26216 16042
rect 25670 7884 25732 9724
rect 26160 7884 26216 9724
rect 35922 14142 36468 14230
rect 35922 12976 35996 14142
rect 36384 12976 36468 14142
rect 33458 9667 34404 9722
rect 33458 8013 33545 9667
rect 34317 8013 34404 9667
rect 33458 7910 34404 8013
rect 25670 7814 26216 7884
rect 98 5787 1136 5814
rect 98 3848 652 5787
rect 1082 3848 1136 5787
rect 35922 5752 36468 12976
rect 44943 9627 46398 9715
rect 44943 8021 45015 9627
rect 46295 8021 46398 9627
rect 44943 7925 46398 8021
rect 27733 5627 28735 5699
rect 25502 5390 25884 5452
rect 25502 4474 25564 5390
rect 25826 4474 25884 5390
rect 25502 4406 25884 4474
rect 27733 4029 27804 5627
rect 28679 4029 28735 5627
rect 27733 3950 28735 4029
rect 98 3814 1136 3848
rect 35922 3912 35984 5752
rect 36412 3912 36468 5752
rect 38097 5627 39751 5699
rect 38097 4021 38176 5627
rect 39679 4021 39751 5627
rect 38097 3942 39751 4021
rect 35922 3830 36468 3912
rect 79605 1360 80693 1539
rect 78651 1003 79232 1004
rect 79605 1003 79784 1360
rect 46343 954 46692 955
rect 46343 807 46344 954
rect 46691 807 76672 954
rect 78651 824 78652 1003
rect 79231 824 79784 1003
rect 78651 823 79232 824
rect 46343 806 46692 807
rect 76525 236 76672 807
rect 76525 89 80685 236
<< via4 >>
rect 9792 23427 10155 23788
rect 26800 22916 27164 23264
rect 29708 23213 30098 23214
rect 29708 22825 29709 23213
rect 29709 22825 30097 23213
rect 30097 22825 30098 23213
rect 29708 22824 30098 22825
rect 40777 23094 41167 23095
rect 40777 22706 40778 23094
rect 40778 22706 41166 23094
rect 41166 22706 41167 23094
rect 40777 22705 41167 22706
rect 82573 22795 83368 23579
rect 82564 22319 83366 22320
rect 82564 21519 82565 22319
rect 82565 21519 83365 22319
rect 83365 21519 83366 22319
rect 82564 21518 83366 21519
rect 6405 17856 6891 19773
rect 82564 19233 83366 19234
rect 26592 18488 26894 18796
rect 31778 18585 32279 18586
rect 31778 18086 31779 18585
rect 31779 18086 32278 18585
rect 32278 18086 32279 18585
rect 31778 18085 32279 18086
rect 43168 18867 43558 18868
rect 43168 18479 43169 18867
rect 43169 18479 43557 18867
rect 43557 18479 43558 18867
rect 43168 18478 43558 18479
rect 82564 18433 82565 19233
rect 82565 18433 83365 19233
rect 83365 18433 83366 19233
rect 82564 18432 83366 18433
rect 846 7841 1276 9780
rect 25734 16042 26134 17396
rect 25732 7884 26160 9724
rect 35996 12976 36384 14142
rect 33545 8013 34317 9667
rect 652 3848 1082 5787
rect 45015 8021 46295 9627
rect 82564 9357 83366 9358
rect 82564 8557 82565 9357
rect 82565 8557 83365 9357
rect 83365 8557 83366 9357
rect 82564 8556 83366 8557
rect 25564 4474 25826 5390
rect 27804 4029 28679 5627
rect 35984 3912 36412 5752
rect 38176 4021 39679 5627
rect 82564 5045 83366 5046
rect 82564 4245 82565 5045
rect 82565 4245 83365 5045
rect 83365 4245 83366 5045
rect 82564 4244 83366 4245
rect 80693 1290 81413 1610
rect 80685 3 81405 323
<< metal5 >>
rect 1 23788 84138 23813
rect 1 23427 9792 23788
rect 10155 23579 84138 23788
rect 10155 23427 82573 23579
rect 1 23264 82573 23427
rect 1 22916 26800 23264
rect 27164 23214 82573 23264
rect 27164 22916 29708 23214
rect 1 22824 29708 22916
rect 30098 23095 82573 23214
rect 30098 22824 40777 23095
rect 1 22705 40777 22824
rect 41167 22795 82573 23095
rect 83368 22795 84138 23579
rect 41167 22705 84138 22795
rect 1 22320 84138 22705
rect 1 21813 82564 22320
rect 82540 21518 82564 21813
rect 83366 21813 84138 22320
rect 83366 21518 83390 21813
rect 82540 21494 83390 21518
rect 1 19773 84138 19813
rect 1 17856 6405 19773
rect 6891 19234 84138 19773
rect 6891 18868 82564 19234
rect 6891 18796 43168 18868
rect 6891 18488 26592 18796
rect 26894 18586 43168 18796
rect 26894 18488 31778 18586
rect 6891 18085 31778 18488
rect 32279 18478 43168 18586
rect 43558 18478 82564 18868
rect 32279 18432 82564 18478
rect 83366 18432 84138 19234
rect 32279 18085 84138 18432
rect 6891 17856 84138 18085
rect 1 17813 84138 17856
rect 25654 17468 26220 17476
rect 25654 17396 47138 17468
rect 25654 16042 25734 17396
rect 26134 17134 47138 17396
rect 26134 16042 26220 17134
rect 25654 15970 26220 16042
rect 27552 15576 46128 16082
rect 35920 14142 36470 15576
rect 35920 12976 35996 14142
rect 36384 12976 36470 14142
rect 35920 12882 36470 12976
rect 1 9780 84186 9813
rect 1 7841 846 9780
rect 1276 9724 84186 9780
rect 1276 7884 25732 9724
rect 26160 9667 84186 9724
rect 26160 8013 33545 9667
rect 34317 9627 84186 9667
rect 34317 8021 45015 9627
rect 46295 9358 84186 9627
rect 46295 8556 82564 9358
rect 83366 8556 84186 9358
rect 46295 8021 84186 8556
rect 34317 8013 84186 8021
rect 26160 7884 84186 8013
rect 1276 7841 84186 7884
rect 1 7813 84186 7841
rect 1 5787 84186 5813
rect 1 3848 652 5787
rect 1082 5752 84186 5787
rect 1082 5627 35984 5752
rect 1082 5390 27804 5627
rect 1082 4474 25564 5390
rect 25826 4474 27804 5390
rect 1082 4029 27804 4474
rect 28679 4029 35984 5627
rect 1082 3912 35984 4029
rect 36412 5627 84186 5752
rect 36412 4021 38176 5627
rect 39679 5046 84186 5627
rect 39679 4244 82564 5046
rect 83366 4244 84186 5046
rect 39679 4021 84186 4244
rect 36412 3912 84186 4021
rect 1082 3848 84186 3912
rect 1 3813 84186 3848
rect 80669 1610 81437 1634
rect 80669 1600 80693 1610
rect 80668 1290 80693 1600
rect 81413 1600 81437 1610
rect 81413 1290 84200 1600
rect 80668 1280 84200 1290
rect 80669 1266 81437 1280
rect 80661 323 81429 347
rect 80661 320 80685 323
rect 80660 3 80685 320
rect 81405 320 81429 323
rect 81405 3 84200 320
rect 80660 0 84200 3
rect 80661 -21 81429 0
use sky130_be_ip__lsxo  sky130_be_ip__lsxo_0 ../ip/sky130_be_ip__lsxo/mag
timestamp 1714591373
transform 1 0 -202 0 1 24278
box 1476 -23704 25570 -812
use sky130_ef_ip__rc_osc_16M  sky130_ef_ip__rc_osc_16M_0 ../ip/sky130_ef_ip__rc_osc_16M/mag
timestamp 1721245376
transform 0 -1 36464 1 0 2774
box 0 700 10977 10024
use sky130_ef_ip__rc_osc_500k  sky130_ef_ip__rc_osc_500k_0 ../ip/sky130_ef_ip__rc_osc_500k/mag
timestamp 1721241604
transform 0 -1 47544 1 0 2698
box 0 0 12242 10724
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_0
array 0 0 2752 0 7 -2622
timestamp 1721093827
transform 0 -1 27659 1 0 16081
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_1
array 0 0 2676 0 6 -2576
timestamp 1721093827
transform 0 -1 31359 1 0 20739
box -1349 -1081 1371 1081
use sky130_ht_ip__hsxo_cpz1  sky130_ht_ip__hsxo_cpz1_0 ../ip/sky130_ht_ip__hsxo_cpz1/mag
timestamp 1718126100
transform -1 0 80215 0 -1 18009
box -3162 -7320 32492 17749
use xres_buf  xres_buf_0
timestamp 1719932489
transform -1 0 29928 0 1 18834
box 284 -400 3656 3800
<< labels >>
flabel metal2 9000 0 9300 300 0 FreeSans 480 90 0 0 lsxo_xin
port 1 nsew
flabel metal2 31000 0 31300 300 0 FreeSans 480 90 0 0 lsxo_xout
port 2 nsew
flabel metal2 53000 0 53300 300 0 FreeSans 480 90 0 0 hsxo_xin
port 3 nsew
flabel metal2 75000 0 75300 300 0 FreeSans 480 90 0 0 hsxo_xout
port 4 nsew
flabel metal2 32400 25300 32428 25600 0 FreeSans 480 90 0 0 rc_osc_16M_ena
port 5 nsew
flabel metal2 32848 25300 32876 25600 0 FreeSans 480 90 0 0 rc_osc_500k_ena
port 6 nsew
flabel metal2 33296 25300 33324 25600 0 FreeSans 480 90 0 0 lsxo_ena
port 7 nsew
flabel metal2 33744 25300 33772 25600 0 FreeSans 480 90 0 0 lsxo_standby
port 8 nsew
flabel metal2 34192 25300 34220 25600 0 FreeSans 480 90 0 0 hsxo_ena
port 9 nsew
flabel metal2 34640 25300 34668 25600 0 FreeSans 480 90 0 0 hsxo_standby
port 10 nsew
flabel metal2 35088 25300 35116 25600 0 FreeSans 480 90 0 0 rc_osc_16M_dout
port 11 nsew
flabel metal2 35536 25300 35564 25600 0 FreeSans 480 90 0 0 rc_osc_500k_dout
port 12 nsew
flabel metal2 35984 25300 36012 25600 0 FreeSans 480 90 0 0 lsxo_dout
port 13 nsew
flabel metal2 36432 25300 36460 25600 0 FreeSans 480 90 0 0 hsxo_dout
port 14 nsew
flabel metal5 83560 0 84200 320 0 FreeSans 800 0 0 0 lsxo_ibias
port 15 nsew
flabel metal5 83560 1280 84200 1600 0 FreeSans 800 0 0 0 hsxo_ibias
port 16 nsew
flabel metal2 31504 25300 31532 25600 0 FreeSans 480 90 0 0 resetb_in_h
port 22 nsew
flabel metal2 31952 25300 31980 25600 0 FreeSans 480 90 0 0 resetb_out_l
port 23 nsew
flabel metal5 83697 3813 84186 5813 0 FreeSans 3200 90 0 0 vdda3
port 19 nsew
flabel metal5 83697 7813 84186 9813 0 FreeSans 3200 90 0 0 vssa3
port 17 nsew
flabel metal5 83649 17813 84138 19813 0 FreeSans 3200 90 0 0 vccd0
port 20 nsew
flabel metal5 83649 21813 84138 23813 0 FreeSans 3200 90 0 0 vssd0
port 21 nsew
flabel metal5 1 3813 652 5813 0 FreeSans 3200 90 0 0 vdda3
port 19 nsew
flabel metal5 1 7813 846 9813 0 FreeSans 3200 90 0 0 vssa3
port 17 nsew
flabel metal5 1 17813 601 19813 0 FreeSans 3200 90 0 0 vccd0
port 20 nsew
flabel metal5 1 21813 601 23813 0 FreeSans 3200 90 0 0 vssd0
port 21 nsew
<< properties >>
string FIXED_BBOX 0 0 84186 25676
<< end >>
