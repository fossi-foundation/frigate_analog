VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_routes_user
  CLASS COVER ;
  FOREIGN analog_routes_user ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 100.000 ;
  OBS
      LAYER met4 ;
        RECT 0.000 2.210 0.640 100.000 ;
        RECT 1.280 0.000 1.920 100.000 ;
        RECT 2.560 2.210 3.200 100.000 ;
        RECT 3.840 0.000 4.480 100.000 ;
        RECT 5.120 2.210 5.760 100.000 ;
        RECT 6.400 0.000 7.040 100.000 ;
        RECT 7.680 2.210 8.320 100.000 ;
        RECT 8.960 0.000 9.600 100.000 ;
        RECT 10.240 2.210 10.880 100.000 ;
        RECT 11.520 0.000 12.160 100.000 ;
        RECT 12.800 2.210 13.440 100.000 ;
        RECT 14.080 0.000 14.720 100.000 ;
        RECT 15.360 2.210 16.000 100.000 ;
        RECT 16.640 0.000 17.280 100.000 ;
        RECT 17.920 2.210 18.560 100.000 ;
        RECT 19.200 0.000 19.840 100.000 ;
        RECT 20.480 2.210 21.120 100.000 ;
        RECT 21.760 0.000 22.400 100.000 ;
        RECT 23.040 2.210 23.680 100.000 ;
        RECT 24.320 0.000 24.960 100.000 ;
        RECT 25.600 2.210 26.240 100.000 ;
        RECT 26.880 0.000 27.520 100.000 ;
        RECT 28.160 2.210 28.800 100.000 ;
        RECT 29.440 0.000 30.080 100.000 ;
        RECT 30.720 2.210 31.360 100.000 ;
        RECT 32.000 0.000 32.640 100.000 ;
        RECT 33.280 2.210 33.920 100.000 ;
        RECT 34.560 0.000 35.200 100.000 ;
        RECT 35.840 2.210 36.480 100.000 ;
        RECT 37.120 0.000 37.760 100.000 ;
        RECT 38.400 2.210 39.040 100.000 ;
        RECT 39.680 0.000 40.320 100.000 ;
        RECT 40.960 2.210 41.600 100.000 ;
        RECT 42.240 0.000 42.880 100.000 ;
        RECT 43.520 2.210 44.160 100.000 ;
        RECT 44.800 0.000 45.440 100.000 ;
        RECT 46.080 2.210 46.720 100.000 ;
        RECT 47.360 0.000 48.000 100.000 ;
        RECT 48.640 2.210 49.280 100.000 ;
        RECT 49.920 0.000 50.560 100.000 ;
        RECT 51.200 2.210 51.840 100.000 ;
        RECT 52.480 0.000 53.120 100.000 ;
        RECT 53.760 2.210 54.400 100.000 ;
        RECT 55.040 0.000 55.680 100.000 ;
        RECT 56.320 2.210 56.960 100.000 ;
        RECT 57.600 0.000 58.240 100.000 ;
        RECT 58.880 2.210 59.520 100.000 ;
        RECT 60.160 0.000 60.800 100.000 ;
        RECT 61.440 2.210 62.080 100.000 ;
        RECT 62.720 0.000 63.360 100.000 ;
        RECT 64.000 2.210 64.640 100.000 ;
        RECT 65.280 0.000 65.920 100.000 ;
        RECT 66.560 2.210 67.200 100.000 ;
        RECT 67.840 0.000 68.480 100.000 ;
        RECT 69.120 2.210 69.760 100.000 ;
        RECT 70.400 0.000 71.040 100.000 ;
        RECT 71.680 2.210 72.320 100.000 ;
        RECT 72.960 0.000 73.600 100.000 ;
        RECT 74.240 2.210 74.880 100.000 ;
        RECT 75.520 0.000 76.160 100.000 ;
        RECT 76.800 2.210 77.440 100.000 ;
        RECT 78.080 0.000 78.720 100.000 ;
        RECT 79.360 2.210 80.000 100.000 ;
  END
END analog_routes_user
END LIBRARY

