magic
tech sky130A
magscale 1 2
timestamp 1724444054
<< metal1 >>
rect -372 11602 -336 23127
rect -288 11729 -252 23127
rect -296 11723 -252 11729
rect -301 11671 -295 11723
rect -243 11671 -237 11723
rect -296 11665 -252 11671
rect -288 11644 -252 11665
rect -382 11596 -336 11602
rect -384 11544 -378 11596
rect -326 11544 -320 11596
rect -382 11538 -336 11544
rect -372 11529 -336 11538
rect -204 5682 -168 23127
rect -120 5809 -84 23127
rect -36 18182 0 23127
rect 48 18309 84 23127
rect 40 18303 84 18309
rect 1008 18673 1208 18680
rect 1008 18466 5616 18673
rect 35 18251 41 18303
rect 93 18251 99 18303
rect 40 18245 84 18251
rect 48 18241 84 18245
rect -46 18176 0 18182
rect -48 18124 -42 18176
rect 10 18124 16 18176
rect -46 18118 0 18124
rect 9 17768 221 17790
rect 9 17363 36 17768
rect 200 17363 221 17768
rect 9 16848 221 17363
rect 18 10942 218 12650
rect 1008 12063 1208 18466
rect 1749 18252 1755 18304
rect 1807 18252 1813 18304
rect 1462 18177 1511 18197
rect 1455 18125 1461 18177
rect 1513 18125 1519 18177
rect 1462 16848 1511 18125
rect 1756 16813 1805 18252
rect 5409 17545 5616 18466
rect 7498 18182 7534 23127
rect 7582 18309 7618 23127
rect 7574 18303 7618 18309
rect 7569 18251 7575 18303
rect 7627 18251 7633 18303
rect 7574 18245 7618 18251
rect 7582 18241 7618 18245
rect 7488 18176 7534 18182
rect 7486 18124 7492 18176
rect 7544 18124 7550 18176
rect 7488 18118 7534 18124
rect 5409 17519 7574 17545
rect 5409 17366 7233 17519
rect 7546 17366 7574 17519
rect 5409 17338 7574 17366
rect 1008 11856 5608 12063
rect -128 5803 -84 5809
rect -133 5751 -127 5803
rect -75 5751 -69 5803
rect -128 5745 -84 5751
rect -120 5741 -84 5745
rect -214 5676 -168 5682
rect -216 5624 -210 5676
rect -158 5624 -152 5676
rect -214 5618 -168 5624
rect 18 5042 218 6728
rect 1008 5848 1208 11856
rect 1756 11724 1805 11753
rect 1749 11672 1755 11724
rect 1807 11672 1813 11724
rect 1462 11597 1511 11619
rect 1455 11545 1461 11597
rect 1513 11545 1519 11597
rect 1462 10926 1511 11545
rect 1756 10913 1805 11672
rect 5401 11448 5608 11856
rect 7666 11602 7702 23127
rect 7750 11729 7786 23127
rect 7742 11723 7786 11729
rect 7737 11671 7743 11723
rect 7795 11671 7801 11723
rect 7742 11665 7786 11671
rect 7750 11644 7786 11665
rect 7656 11596 7702 11602
rect 7654 11544 7660 11596
rect 7712 11544 7718 11596
rect 7656 11538 7702 11544
rect 7666 11529 7702 11538
rect 7210 11448 7762 11450
rect 5401 11422 7762 11448
rect 5401 11255 7239 11422
rect 7726 11255 7762 11422
rect 5401 11241 7762 11255
rect 7210 11235 7762 11241
rect 1008 5579 1214 5848
rect 1756 5804 1805 5824
rect 1749 5752 1755 5804
rect 1807 5752 1813 5804
rect 1462 5677 1511 5695
rect 1455 5625 1461 5677
rect 1513 5625 1519 5677
rect 1008 6 1208 5579
rect 1462 5004 1511 5625
rect 1756 5004 1805 5752
rect 7834 5682 7870 23127
rect 7918 5809 7954 23127
rect 8032 18395 8232 23148
rect 9082 18395 9246 23151
rect 9506 23066 9576 23134
rect 9800 23066 9870 23134
rect 8032 18066 8262 18395
rect 9082 18255 9256 18395
rect 8032 16200 8232 18066
rect 9052 17956 9256 18255
rect 9787 18252 9793 18304
rect 9845 18252 9851 18304
rect 9500 18177 9549 18197
rect 9493 18125 9499 18177
rect 9551 18125 9557 18177
rect 9046 17539 9256 17956
rect 9042 17507 9256 17539
rect 9042 17052 9068 17507
rect 9045 16852 9068 17052
rect 9046 16756 9068 16852
rect 9226 16756 9246 17507
rect 9500 16848 9549 18125
rect 9794 16813 9843 18252
rect 8056 10960 8256 12631
rect 9046 11393 9246 16756
rect 9794 11724 9843 11733
rect 9787 11672 9793 11724
rect 9845 11672 9851 11724
rect 9500 11597 9549 11606
rect 9493 11545 9499 11597
rect 9551 11545 9557 11597
rect 9046 11353 9271 11393
rect 9046 10766 9084 11353
rect 9252 10766 9271 11353
rect 9500 10926 9549 11545
rect 9794 10913 9843 11672
rect 15704 11602 15740 23127
rect 15788 11729 15824 23127
rect 15780 11723 15824 11729
rect 15775 11671 15781 11723
rect 15833 11671 15839 11723
rect 15780 11665 15824 11671
rect 15788 11663 15824 11665
rect 15694 11596 15740 11602
rect 15692 11544 15698 11596
rect 15750 11544 15756 11596
rect 15694 11538 15740 11544
rect 15704 11537 15740 11538
rect 9046 10732 9271 10766
rect 7910 5803 7954 5809
rect 7905 5751 7911 5803
rect 7963 5751 7969 5803
rect 7910 5745 7954 5751
rect 7918 5741 7954 5745
rect 7824 5676 7870 5682
rect 7822 5624 7828 5676
rect 7880 5624 7886 5676
rect 7824 5618 7870 5624
rect 8056 5078 8256 6728
rect 9046 5848 9246 10732
rect 9046 5579 9252 5848
rect 9794 5804 9843 5824
rect 9787 5752 9793 5804
rect 9845 5752 9851 5804
rect 9500 5677 9549 5695
rect 9493 5625 9499 5677
rect 9551 5625 9557 5677
rect 9046 6 9246 5579
rect 9500 5004 9549 5625
rect 9794 5004 9843 5752
rect 15872 5682 15908 23127
rect 15956 5809 15992 23127
rect 16040 18182 16076 23127
rect 16124 18309 16160 23127
rect 16116 18303 16160 18309
rect 16111 18251 16117 18303
rect 16169 18251 16175 18303
rect 17825 18252 17831 18304
rect 17883 18252 17889 18304
rect 16116 18245 16160 18251
rect 16124 18241 16160 18245
rect 16030 18176 16076 18182
rect 17538 18177 17587 18197
rect 16028 18124 16034 18176
rect 16086 18124 16092 18176
rect 17531 18125 17537 18177
rect 17589 18125 17595 18177
rect 16030 18118 16076 18124
rect 17538 16848 17587 18125
rect 17832 16813 17881 18252
rect 23574 18182 23610 23127
rect 23658 18309 23694 23127
rect 23650 18303 23694 18309
rect 23645 18251 23651 18303
rect 23703 18251 23709 18303
rect 23650 18245 23694 18251
rect 23658 18241 23694 18245
rect 23564 18176 23610 18182
rect 23562 18124 23568 18176
rect 23620 18124 23626 18176
rect 23564 18118 23610 18124
rect 16108 16304 16122 16628
rect 16094 11004 16294 12650
rect 17084 11447 17284 16664
rect 17832 11724 17881 11733
rect 17825 11672 17831 11724
rect 17883 11672 17889 11724
rect 17538 11597 17587 11602
rect 17531 11545 17537 11597
rect 17589 11545 17595 11597
rect 17090 11393 17284 11447
rect 17090 11353 17299 11393
rect 17090 10766 17112 11353
rect 17280 10766 17299 11353
rect 17538 10926 17587 11545
rect 17832 10913 17881 11672
rect 23742 11602 23778 23127
rect 23826 11729 23862 23127
rect 23818 11723 23862 11729
rect 23813 11671 23819 11723
rect 23871 11671 23877 11723
rect 23818 11665 23862 11671
rect 23826 11644 23862 11665
rect 23732 11596 23778 11602
rect 23730 11544 23736 11596
rect 23788 11544 23794 11596
rect 23732 11538 23778 11544
rect 23742 11529 23778 11538
rect 17090 10732 17299 10766
rect 17090 10713 17284 10732
rect 15948 5803 15992 5809
rect 15943 5751 15949 5803
rect 16001 5751 16007 5803
rect 15948 5745 15992 5751
rect 15956 5741 15992 5745
rect 15862 5676 15908 5682
rect 15860 5624 15866 5676
rect 15918 5624 15924 5676
rect 15862 5618 15908 5624
rect 16094 5060 16294 6728
rect 17084 5848 17284 10713
rect 17084 5579 17290 5848
rect 17832 5804 17881 5824
rect 17825 5752 17831 5804
rect 17883 5752 17889 5804
rect 17538 5677 17587 5695
rect 17531 5625 17537 5677
rect 17589 5625 17595 5677
rect 17084 6 17284 5579
rect 17538 5004 17587 5625
rect 17832 5004 17881 5752
rect 23910 5682 23946 23127
rect 23994 5809 24030 23127
rect 24138 16922 24338 18746
rect 25128 14236 25328 23137
rect 25568 23072 25638 23140
rect 25860 23070 25930 23138
rect 25863 18252 25869 18304
rect 25921 18252 25927 18304
rect 25576 18177 25625 18197
rect 25569 18125 25575 18177
rect 25627 18125 25633 18177
rect 25576 17023 25625 18125
rect 25870 16813 25919 18252
rect 25128 14218 25334 14236
rect 25128 13422 25153 14218
rect 25314 13422 25334 14218
rect 25128 13405 25334 13422
rect 24132 10978 24332 12650
rect 23986 5803 24030 5809
rect 23981 5751 23987 5803
rect 24039 5751 24045 5803
rect 23986 5745 24030 5751
rect 23994 5741 24030 5745
rect 23900 5676 23946 5682
rect 23898 5624 23904 5676
rect 23956 5624 23962 5676
rect 23900 5618 23946 5624
rect 24132 5076 24332 6728
rect 25128 6 25328 13405
rect 25870 11724 25919 11753
rect 25863 11672 25869 11724
rect 25921 11672 25927 11724
rect 25576 11597 25625 11619
rect 25569 11545 25575 11597
rect 25627 11545 25633 11597
rect 25576 10948 25625 11545
rect 25870 10913 25919 11672
rect 25870 5804 25919 5824
rect 25863 5752 25869 5804
rect 25921 5752 25927 5804
rect 25576 5677 25625 5695
rect 25569 5625 25575 5677
rect 25627 5625 25633 5677
rect 25576 5048 25625 5625
rect 25870 5013 25919 5752
<< via1 >>
rect -295 11671 -243 11723
rect -378 11544 -326 11596
rect 41 18251 93 18303
rect -42 18124 10 18176
rect 36 17363 200 17768
rect 1755 18252 1807 18304
rect 1461 18125 1513 18177
rect 7575 18251 7627 18303
rect 7492 18124 7544 18176
rect 7233 17366 7546 17519
rect -127 5751 -75 5803
rect -210 5624 -158 5676
rect 1755 11672 1807 11724
rect 1461 11545 1513 11597
rect 7743 11671 7795 11723
rect 7660 11544 7712 11596
rect 7239 11255 7726 11422
rect 1755 5752 1807 5804
rect 1461 5625 1513 5677
rect 9793 18252 9845 18304
rect 9499 18125 9551 18177
rect 9068 16756 9226 17507
rect 9793 11672 9845 11724
rect 9499 11545 9551 11597
rect 9084 10766 9252 11353
rect 15781 11671 15833 11723
rect 15698 11544 15750 11596
rect 7911 5751 7963 5803
rect 7828 5624 7880 5676
rect 9793 5752 9845 5804
rect 9499 5625 9551 5677
rect 16117 18251 16169 18303
rect 17831 18252 17883 18304
rect 16034 18124 16086 18176
rect 17537 18125 17589 18177
rect 23651 18251 23703 18303
rect 23568 18124 23620 18176
rect 17831 11672 17883 11724
rect 17537 11545 17589 11597
rect 17112 10766 17280 11353
rect 23819 11671 23871 11723
rect 23736 11544 23788 11596
rect 15949 5751 16001 5803
rect 15866 5624 15918 5676
rect 17831 5752 17883 5804
rect 17537 5625 17589 5677
rect 25869 18252 25921 18304
rect 25575 18125 25627 18177
rect 25153 13422 25314 14218
rect 23987 5751 24039 5803
rect 23904 5624 23956 5676
rect 25869 11672 25921 11724
rect 25575 11545 25627 11597
rect 25869 5752 25921 5804
rect 25575 5625 25627 5677
<< metal2 >>
rect 8038 19768 8236 19813
rect 8038 18744 8076 19768
rect 5416 18574 8076 18744
rect 8204 18744 8236 19768
rect 8204 18574 8243 18744
rect 5416 18551 8243 18574
rect 41 18303 93 18309
rect 34 18253 41 18302
rect 1755 18304 1807 18310
rect 93 18253 1755 18302
rect 41 18245 93 18251
rect 1755 18246 1807 18252
rect -42 18176 10 18182
rect -48 18126 -42 18175
rect 1461 18177 1513 18183
rect 10 18126 1461 18175
rect -42 18118 10 18124
rect 1461 18119 1513 18125
rect 5416 17797 5609 18551
rect 8038 18536 8236 18551
rect 7575 18303 7627 18309
rect 9793 18304 9845 18310
rect 7627 18253 9793 18302
rect 7575 18245 7627 18251
rect 16117 18303 16169 18309
rect 16113 18253 16117 18302
rect 9793 18246 9845 18252
rect 17831 18304 17883 18310
rect 16169 18253 17831 18302
rect 16117 18245 16169 18251
rect 17831 18246 17883 18252
rect 23651 18303 23703 18309
rect 25869 18304 25921 18310
rect 23703 18253 25869 18302
rect 23651 18245 23703 18251
rect 25869 18246 25921 18252
rect 7492 18176 7544 18182
rect 9499 18177 9551 18183
rect 7544 18126 9499 18175
rect 7492 18118 7544 18124
rect 16034 18176 16086 18182
rect 16027 18126 16034 18175
rect 9499 18119 9551 18125
rect 17537 18177 17589 18183
rect 16086 18126 17537 18175
rect 16034 18118 16086 18124
rect 17537 18119 17589 18125
rect 23568 18176 23620 18182
rect 25575 18177 25627 18183
rect 23620 18126 25575 18175
rect 23568 18118 23620 18124
rect 25575 18119 25627 18125
rect 8 17768 5609 17797
rect 8 17363 36 17768
rect 200 17363 5609 17768
rect 8 17327 5609 17363
rect 6120 17728 31739 17974
rect 8 17322 5605 17327
rect 6120 16666 7093 17728
rect 7206 17519 9257 17542
rect 7206 17366 7233 17519
rect 7546 17507 9257 17519
rect 7546 17366 9068 17507
rect 7206 17342 9068 17366
rect 9042 16756 9068 17342
rect 9226 17342 9257 17507
rect 9226 16756 9246 17342
rect 9042 16731 9246 16756
rect 14158 16662 15131 17728
rect 22196 17128 31717 17374
rect 22196 16638 23169 17128
rect 30234 16666 31207 17128
rect 25133 14218 25334 14236
rect 16072 13481 16299 13516
rect 16072 12497 16102 13481
rect 16276 12497 16299 13481
rect 16072 12463 16299 12497
rect 24079 13450 24298 13493
rect 24079 12487 24112 13450
rect 24258 12487 24298 13450
rect 25133 13422 25153 14218
rect 25314 13422 25334 14218
rect 25133 13405 25334 13422
rect 24079 12448 24298 12487
rect 6120 11806 31739 12052
rect -295 11723 -243 11729
rect 1755 11724 1807 11730
rect -243 11673 1755 11722
rect -295 11665 -243 11671
rect 1755 11666 1807 11672
rect -378 11596 -326 11602
rect 1461 11597 1513 11603
rect -326 11546 1461 11595
rect -378 11538 -326 11544
rect 1461 11539 1513 11545
rect 6120 10744 7093 11806
rect 7743 11723 7795 11729
rect 9793 11724 9845 11730
rect 7795 11673 9793 11722
rect 7743 11665 7795 11671
rect 9793 11666 9845 11672
rect 7660 11596 7712 11602
rect 9499 11597 9551 11603
rect 7712 11546 9499 11595
rect 7660 11538 7712 11544
rect 9499 11539 9551 11545
rect 7210 11422 7762 11450
rect 7210 11255 7239 11422
rect 7726 11417 7762 11422
rect 7726 11353 9274 11417
rect 7726 11255 9084 11353
rect 7210 11241 9084 11255
rect 7210 11235 7762 11241
rect 9050 10766 9084 11241
rect 9252 11241 9274 11353
rect 9252 10766 9271 11241
rect 9050 10732 9271 10766
rect 14158 10742 15131 11806
rect 15781 11723 15833 11729
rect 17831 11724 17883 11730
rect 15833 11673 17831 11722
rect 15781 11665 15833 11671
rect 17831 11666 17883 11672
rect 23819 11723 23871 11729
rect 25869 11724 25921 11730
rect 23871 11673 25869 11722
rect 23819 11665 23871 11671
rect 25869 11666 25921 11672
rect 15698 11596 15750 11602
rect 17537 11597 17589 11603
rect 15750 11546 17537 11595
rect 15698 11538 15750 11544
rect 17537 11539 17589 11545
rect 23736 11596 23788 11602
rect 25575 11597 25627 11603
rect 23788 11546 25575 11595
rect 23736 11538 23788 11544
rect 25575 11539 25627 11545
rect 17083 11353 17299 11393
rect 17083 10766 17112 11353
rect 17280 10766 17299 11353
rect 22156 11206 31759 11452
rect 17083 10732 17299 10766
rect 22196 10740 23169 11206
rect 30234 10742 31207 11206
rect 6120 5884 31801 6130
rect -127 5803 -75 5809
rect 1755 5804 1807 5810
rect -75 5753 1755 5802
rect -127 5745 -75 5751
rect 1755 5746 1807 5752
rect -210 5676 -158 5682
rect 1461 5677 1513 5683
rect -158 5626 1461 5675
rect -210 5618 -158 5624
rect 1461 5619 1513 5625
rect 6120 4766 7093 5884
rect 7911 5803 7963 5809
rect 9793 5804 9845 5810
rect 7963 5753 9793 5802
rect 7911 5745 7963 5751
rect 9793 5746 9845 5752
rect 7828 5676 7880 5682
rect 9499 5677 9551 5683
rect 7880 5626 9499 5675
rect 7828 5618 7880 5624
rect 9499 5619 9551 5625
rect 14158 4818 15131 5884
rect 15949 5803 16001 5809
rect 17831 5804 17883 5810
rect 16001 5753 17831 5802
rect 15949 5745 16001 5751
rect 17831 5746 17883 5752
rect 23987 5803 24039 5809
rect 25869 5804 25921 5810
rect 24039 5753 25869 5802
rect 23987 5745 24039 5751
rect 25869 5746 25921 5752
rect 15866 5676 15918 5682
rect 17537 5677 17589 5683
rect 15918 5626 17537 5675
rect 15866 5618 15918 5624
rect 17537 5619 17589 5625
rect 23904 5676 23956 5682
rect 25575 5677 25627 5683
rect 23956 5626 25575 5675
rect 23904 5618 23956 5624
rect 25575 5619 25627 5625
rect 22184 5272 31779 5518
rect 22196 4814 23169 5272
rect 30234 4812 31207 5272
rect 24071 1562 24305 1590
rect 8019 1458 8248 1490
rect 8019 655 8040 1458
rect 8217 655 8248 1458
rect 8019 628 8248 655
rect 24071 643 24104 1562
rect 24281 643 24305 1562
rect 24071 611 24305 643
<< via2 >>
rect 8076 18574 8204 19768
rect 9068 16756 9226 17507
rect 16102 12497 16276 13481
rect 24112 12487 24258 13450
rect 25153 13422 25314 14218
rect 9084 10766 9252 11353
rect 17112 10766 17280 11353
rect 8040 655 8217 1458
rect 24104 643 24281 1562
<< metal3 >>
rect 8014 19768 8249 23215
rect 7210 18571 7410 18593
rect 7210 18094 7222 18571
rect 7392 18094 7410 18571
rect 2346 17443 2546 17476
rect 2346 16991 2364 17443
rect 2518 16991 2546 17443
rect 2346 4 2546 16991
rect 2668 384 3640 16674
rect 7210 4 7410 18094
rect 8014 18574 8076 19768
rect 8204 18574 8249 19768
rect 8014 11451 8249 18574
rect 8014 11021 8049 11451
rect 8223 11021 8249 11451
rect 8014 1458 8249 11021
rect 8014 655 8040 1458
rect 8217 655 8249 1458
rect 8014 548 8249 655
rect 9040 17507 9281 23177
rect 14164 23046 15136 23098
rect 9040 16756 9068 17507
rect 9226 16756 9281 17507
rect 9040 12484 9281 16756
rect 9040 12054 9067 12484
rect 9241 12054 9281 12484
rect 9040 11353 9281 12054
rect 9040 10766 9084 11353
rect 9252 10766 9281 11353
rect 9040 1 9281 10766
rect 10384 17453 10584 22624
rect 10384 16976 10399 17453
rect 10569 16976 10584 17453
rect 10384 4 10584 16976
rect 10728 16674 11700 23034
rect 10706 16014 11700 16674
rect 15248 18565 15448 22534
rect 15248 18092 15265 18565
rect 15433 18092 15448 18565
rect 10706 392 11678 16014
rect 15248 0 15448 18092
rect 23300 18568 23500 18604
rect 23300 18102 23326 18568
rect 23481 18102 23500 18568
rect 16069 13481 16304 17591
rect 16069 12497 16102 13481
rect 16276 12497 16304 13481
rect 16069 11458 16304 12497
rect 16069 11028 16099 11458
rect 16273 11028 16304 11458
rect 17074 12455 17315 17591
rect 17074 12025 17103 12455
rect 17277 12025 17315 12455
rect 17074 11441 17315 12025
rect 16069 530 16304 11028
rect 17083 11353 17315 11441
rect 17083 10766 17112 11353
rect 17280 10766 17315 11353
rect 17083 10706 17315 10766
rect 17074 33 17315 10706
rect 18436 17450 18636 17473
rect 18436 16984 18459 17450
rect 18614 16984 18636 17450
rect 18436 86 18636 16984
rect 18758 384 19730 16674
rect 23300 34 23500 18102
rect 24073 13450 24308 23174
rect 25135 14236 25376 23209
rect 26788 22770 27758 23062
rect 30210 23042 31182 23096
rect 24073 12487 24112 13450
rect 24258 12487 24308 13450
rect 25133 14218 25376 14236
rect 25133 13422 25153 14218
rect 25314 13422 25376 14218
rect 25133 13405 25376 13422
rect 24073 11466 24308 12487
rect 24073 11036 24120 11466
rect 24294 11036 24308 11466
rect 24073 1562 24308 11036
rect 24073 643 24104 1562
rect 24281 643 24308 1562
rect 24073 507 24308 643
rect 25135 12471 25376 13405
rect 25135 12041 25159 12471
rect 25333 12041 25376 12471
rect 25135 33 25376 12041
rect 26466 17453 26666 22522
rect 26466 16976 26478 17453
rect 26648 16976 26666 17453
rect 26466 0 26666 16976
rect 26788 526 27760 22770
rect 31330 18568 31530 22528
rect 31330 18095 31347 18568
rect 31515 18095 31530 18568
rect 31330 0 31530 18095
<< via3 >>
rect 7222 18094 7392 18571
rect 2364 16991 2518 17443
rect 8049 11021 8223 11451
rect 9067 12054 9241 12484
rect 10399 16976 10569 17453
rect 15265 18092 15433 18565
rect 23326 18102 23481 18568
rect 16099 11028 16273 11458
rect 17103 12025 17277 12455
rect 18459 16984 18614 17450
rect 24120 11036 24294 11466
rect 25159 12041 25333 12471
rect 26478 16976 26648 17453
rect 31347 18095 31515 18568
<< metal4 >>
rect -405 18571 31657 18587
rect -405 18094 7222 18571
rect 7392 18568 31657 18571
rect 7392 18565 23326 18568
rect 7392 18094 15265 18565
rect -405 18092 15265 18094
rect 15433 18102 23326 18565
rect 23481 18102 31347 18568
rect 15433 18095 31347 18102
rect 31515 18095 31657 18568
rect 15433 18092 31657 18095
rect -405 18080 31657 18092
rect -405 17453 31657 17465
rect -405 17443 10399 17453
rect -405 16991 2364 17443
rect 2518 16991 10399 17443
rect -405 16976 10399 16991
rect 10569 17450 26478 17453
rect 10569 16984 18459 17450
rect 18614 16984 26478 17450
rect 10569 16976 26478 16984
rect 26648 16976 31657 17453
rect -405 16958 31657 16976
rect -368 12484 31694 12508
rect -368 12054 9067 12484
rect 9241 12471 31694 12484
rect 9241 12455 25159 12471
rect 9241 12054 17103 12455
rect -368 12025 17103 12054
rect 17277 12041 25159 12455
rect 25333 12041 31694 12471
rect 17277 12025 31694 12041
rect -368 12001 31694 12025
rect -368 11466 31694 11494
rect -368 11458 24120 11466
rect -368 11451 16099 11458
rect -368 11021 8049 11451
rect 8223 11028 16099 11451
rect 16273 11036 24120 11458
rect 24294 11036 31694 11466
rect 16273 11028 31694 11036
rect 8223 11021 31694 11028
rect -368 10987 31694 11021
use cv3_via2_8cut  cv3_via2_8cut_0
timestamp 1719106786
transform 1 0 -4464 0 1 -58458
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_1
timestamp 1719106786
transform 1 0 -4488 0 1 -61482
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_2
timestamp 1719106786
transform 1 0 396 0 1 -58452
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_3
timestamp 1719106786
transform 1 0 402 0 1 -61486
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_4
timestamp 1719106786
transform 1 0 3550 0 1 -61482
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_5
timestamp 1719106786
transform 1 0 3574 0 1 -58458
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_6
timestamp 1719106786
transform 1 0 8440 0 1 -61486
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_7
timestamp 1719106786
transform 1 0 8434 0 1 -58452
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_8
timestamp 1719106786
transform 1 0 11588 0 1 -61482
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_9
timestamp 1719106786
transform 1 0 11612 0 1 -58458
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_10
timestamp 1719106786
transform 1 0 16478 0 1 -61486
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_11
timestamp 1719106786
transform 1 0 16472 0 1 -58452
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_12
timestamp 1719106786
transform 1 0 -4488 0 1 -55560
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_13
timestamp 1719106786
transform 1 0 -4464 0 1 -52536
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_14
timestamp 1719106786
transform 1 0 402 0 1 -55564
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_15
timestamp 1719106786
transform 1 0 396 0 1 -52530
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_16
timestamp 1719106786
transform 1 0 19626 0 1 -61482
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_17
timestamp 1719106786
transform 1 0 19650 0 1 -58458
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_18
timestamp 1719106786
transform 1 0 24516 0 1 -61486
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_19
timestamp 1719106786
transform 1 0 24510 0 1 -58452
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_20
timestamp 1719106786
transform 1 0 19626 0 1 -55560
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_21
timestamp 1719106786
transform 1 0 19650 0 1 -52536
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_22
timestamp 1719106786
transform 1 0 24516 0 1 -55564
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_23
timestamp 1719106786
transform 1 0 24510 0 1 -52530
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_24
timestamp 1719106786
transform 1 0 11588 0 1 -55560
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_25
timestamp 1719106786
transform 1 0 11612 0 1 -52536
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_26
timestamp 1719106786
transform 1 0 16478 0 1 -55564
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_27
timestamp 1719106786
transform 1 0 16472 0 1 -52530
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_28
timestamp 1719106786
transform 1 0 3550 0 1 -55560
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_29
timestamp 1719106786
transform 1 0 3574 0 1 -52536
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_30
timestamp 1719106786
transform 1 0 8440 0 1 -55564
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_31
timestamp 1719106786
transform 1 0 8434 0 1 -52530
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_32
timestamp 1719106786
transform 1 0 3550 0 1 -49638
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_33
timestamp 1719106786
transform 1 0 8440 0 1 -49642
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_34
timestamp 1719106786
transform 1 0 8434 0 1 -46608
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_35
timestamp 1719106786
transform 1 0 3574 0 1 -46614
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_36
timestamp 1719106786
transform 1 0 -4464 0 1 -46614
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_37
timestamp 1719106786
transform 1 0 396 0 1 -46608
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_38
timestamp 1719106786
transform 1 0 402 0 1 -49642
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_39
timestamp 1719106786
transform 1 0 -4488 0 1 -49638
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_40
timestamp 1719106786
transform 1 0 19626 0 1 -49638
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_41
timestamp 1719106786
transform 1 0 16478 0 1 -49642
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_42
timestamp 1719106786
transform 1 0 16472 0 1 -46608
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_43
timestamp 1719106786
transform 1 0 19650 0 1 -46614
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_44
timestamp 1719106786
transform 1 0 11588 0 1 -49638
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_45
timestamp 1719106786
transform 1 0 11612 0 1 -46614
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_46
timestamp 1719106786
transform 1 0 24516 0 1 -49642
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_47
timestamp 1719106786
transform 1 0 24510 0 1 -46608
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_48
timestamp 1719106786
transform 1 0 3558 0 1 -43716
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_49
timestamp 1719106786
transform 1 0 8448 0 1 -43720
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_50
timestamp 1719106786
transform 1 0 3582 0 1 -40692
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_51
timestamp 1719106786
transform 1 0 8442 0 1 -40686
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_52
timestamp 1719106786
transform 1 0 19626 0 1 -43716
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_53
timestamp 1719106786
transform 1 0 24516 0 1 -43720
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_54
timestamp 1719106786
transform 1 0 19650 0 1 -40692
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_55
timestamp 1719106786
transform 1 0 24510 0 1 -40686
box 6850 62208 6998 62544
use cv3_via2_36cut  cv3_via2_36cut_0
timestamp 1719173892
transform 1 0 -544550 0 1 -81734
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_1
timestamp 1719173892
transform 1 0 -552588 0 1 -87694
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_2
timestamp 1719173892
transform 1 0 -544550 0 1 -87662
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_3
timestamp 1719173892
transform 1 0 -536513 0 1 -87671
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_4
timestamp 1719173892
transform 1 0 -528482 0 1 -87694
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_5
timestamp 1719173892
transform 1 0 -528492 0 1 -81778
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_6
timestamp 1719173892
transform 1 0 -536515 0 1 -81776
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_7
timestamp 1719173892
transform 1 0 -536513 0 1 -75861
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_8
timestamp 1719173892
transform 1 0 -528492 0 1 -75860
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_9
timestamp 1719173892
transform 1 0 -528472 0 1 -69744
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_10
timestamp 1719173892
transform 1 0 -544520 0 1 -69714
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_11
timestamp 1719173892
transform 1 0 -552589 0 1 -81766
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_12
timestamp 1719173892
transform 1 0 -541092 0 1 -69456
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_13
timestamp 1719173892
transform 1 0 -544550 0 1 -75850
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_14
timestamp 1719173892
transform 1 0 -552586 0 1 -75836
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_15
timestamp 1719173892
transform 1 0 -525046 0 1 -69456
box 555256 92202 556228 92502
use isolated_switch_xlarge  isolated_switch_xlarge_0 ../ip/sky130_ef_ip__analog_switches/mag
array 0 0 4826 0 1 -16060
timestamp 1724442184
transform 0 -1 9396 -1 0 23810
box 660 -6310 5544 1338
use isolated_switch_xlarge  isolated_switch_xlarge_1
array 0 2 5922 0 3 -8038
timestamp 1724442184
transform 0 -1 1336 -1 0 17714
box 660 -6310 5544 1338
<< labels >>
flabel metal1 17090 10930 17112 11130 0 FreeSans 256 90 0 0 dvdd
port 5 nsew
flabel metal3 11154 17608 11154 17608 0 FreeSans 960 90 0 0 analog1_core
flabel metal3 27258 17608 27258 17608 0 FreeSans 960 90 0 0 analog0_core
flabel metal4 2354 18308 2354 18308 0 FreeSans 1600 0 0 0 avss
flabel metal4 3166 17204 3166 17204 0 FreeSans 1600 0 0 0 avdd
flabel metal4 510 12212 510 12212 0 FreeSans 1600 0 0 0 dvdd
flabel metal4 510 11224 510 11224 0 FreeSans 1600 0 0 0 dvss
flabel metal3 3198 5836 3198 5836 0 FreeSans 960 90 0 0 amuxbusB
flabel metal3 19214 5588 19214 5588 0 FreeSans 960 90 0 0 amuxbusA
flabel metal3 14618 23078 14618 23078 0 FreeSans 960 0 0 0 analog1
flabel metal3 30654 23076 30654 23076 0 FreeSans 960 0 0 0 analog0
flabel metal1 25594 23108 25594 23108 0 FreeSans 480 90 0 0 analog0_connect[1]
flabel metal1 25892 23110 25892 23110 0 FreeSans 480 90 0 0 analog0_connect[0]
flabel metal1 9836 23102 9836 23102 0 FreeSans 480 90 0 0 analog1_connect[0]
flabel metal1 9538 23104 9538 23104 0 FreeSans 480 90 0 0 analog1_connect[1]
flabel metal2 28926 5410 28926 5410 0 FreeSans 960 0 0 0 left_lp_opamp_out
flabel metal2 28882 5988 28882 5988 0 FreeSans 960 0 0 0 left_instramp_out
flabel metal2 28968 11332 28968 11332 0 FreeSans 960 0 0 0 right_hgbw_opamp_out
flabel metal2 29078 11916 29078 11916 0 FreeSans 960 0 0 0 left_hgbw_opamp_out
flabel metal2 29048 17250 29048 17250 0 FreeSans 960 0 0 0 right_instramp_out
flabel metal2 29008 17854 29008 17854 0 FreeSans 960 0 0 0 right_lp_opamp_out
<< end >>
