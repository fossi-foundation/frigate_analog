magic
tech sky130A
magscale 1 2
timestamp 1717861592
<< checkpaint >>
rect -1122 31869 2114 32428
rect -1366 31850 3222 31869
rect -1379 -371 3452 31850
rect -1260 -1260 3060 -371
<< metal2 >>
rect 131 30949 493 30969
rect 131 30655 157 30949
rect 466 30655 493 30949
rect 131 30630 493 30655
rect 749 30947 1400 30969
rect 749 30653 960 30947
rect 1269 30653 1400 30947
rect 749 30630 1400 30653
<< via2 >>
rect 157 30655 466 30949
rect 960 30653 1269 30947
<< metal3 >>
rect 131 30949 600 30969
rect 131 30946 157 30949
rect 466 30946 600 30949
rect 131 30655 155 30946
rect 569 30655 600 30946
rect 131 30630 600 30655
rect 931 30947 1400 30969
rect 931 30656 958 30947
rect 1372 30656 1400 30947
rect 931 30653 960 30656
rect 1269 30653 1400 30656
rect 931 30630 1400 30653
<< via3 >>
rect 155 30655 157 30946
rect 157 30655 466 30946
rect 466 30655 569 30946
rect 958 30656 960 30947
rect 960 30656 1269 30947
rect 1269 30656 1372 30947
<< metal4 >>
rect 131 30946 600 30969
rect 131 30655 155 30946
rect 569 30655 600 30946
rect 131 30630 600 30655
rect 931 30947 1400 30969
rect 931 30656 958 30947
rect 1372 30656 1400 30947
rect 931 30630 1400 30656
rect 0 0 200 30446
rect 400 0 600 30630
rect 800 0 1000 30446
rect 1200 0 1400 30630
rect 1600 0 1800 30446
<< properties >>
string FIXED_BBOX 0 0 1800 30969
string LEFclass COVER
<< end >>
