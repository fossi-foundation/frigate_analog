VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_routes_bottom
  CLASS COVER ;
  FOREIGN analog_routes_bottom ;
  ORIGIN 0.000 0.000 ;
  SIZE 1510.590 BY 112.900 ;
  OBS
      LAYER met2 ;
        RECT 1226.265 53.710 1227.570 55.680 ;
        RECT 1228.430 53.705 1229.735 55.675 ;
        RECT 1273.350 53.625 1274.655 55.595 ;
        RECT 1389.845 53.110 1391.180 55.210 ;
      LAYER met3 ;
        RECT 1226.265 53.710 1227.570 55.680 ;
        RECT 1228.430 53.705 1229.735 55.675 ;
        RECT 1273.350 53.625 1274.655 55.595 ;
        RECT 1389.305 53.105 1391.180 56.175 ;
      LAYER met4 ;
        RECT 1190.075 112.665 1193.275 112.780 ;
        RECT 1190.040 111.180 1193.275 112.665 ;
        RECT 1190.040 15.560 1191.640 111.180 ;
        RECT 1193.310 107.680 1195.210 107.860 ;
        RECT 1193.310 106.080 1196.630 107.680 ;
        RECT 1193.310 105.960 1195.210 106.080 ;
        RECT 1188.480 13.960 1191.680 15.560 ;
        RECT 1193.540 12.205 1195.140 105.960 ;
        RECT 1197.135 102.310 1200.335 102.795 ;
        RECT 1197.040 101.195 1200.335 102.310 ;
        RECT 1193.395 12.055 1195.295 12.205 ;
        RECT 1191.905 10.455 1195.295 12.055 ;
        RECT 1193.395 10.305 1195.295 10.455 ;
        RECT 1197.040 8.610 1198.640 101.195 ;
        RECT 1200.390 97.720 1202.290 97.900 ;
        RECT 1200.390 96.120 1203.710 97.720 ;
        RECT 1200.390 96.000 1202.290 96.120 ;
        RECT 1195.415 7.155 1198.640 8.610 ;
        RECT 1195.415 7.010 1198.615 7.155 ;
        RECT 1200.540 5.235 1202.140 96.000 ;
        RECT 1204.040 92.740 1205.640 93.120 ;
        RECT 1204.040 91.140 1207.365 92.740 ;
        RECT 1200.295 5.165 1202.195 5.235 ;
        RECT 1198.840 3.565 1202.195 5.165 ;
        RECT 1200.295 3.335 1202.195 3.565 ;
        RECT 1204.040 1.720 1205.640 91.140 ;
        RECT 1226.040 87.890 1227.820 87.895 ;
        RECT 1225.985 87.710 1227.885 87.890 ;
        RECT 1225.985 86.110 1229.305 87.710 ;
        RECT 1225.985 85.990 1227.885 86.110 ;
        RECT 1226.205 53.655 1227.630 85.990 ;
        RECT 1228.140 77.740 1230.040 77.920 ;
        RECT 1228.140 76.140 1231.460 77.740 ;
        RECT 1228.140 76.020 1230.040 76.140 ;
        RECT 1228.335 53.615 1229.780 76.020 ;
        RECT 1273.040 67.705 1274.940 67.885 ;
        RECT 1273.040 66.105 1276.360 67.705 ;
        RECT 1273.040 65.985 1274.940 66.105 ;
        RECT 1273.255 53.540 1274.755 65.985 ;
        RECT 1389.310 57.845 1391.180 58.015 ;
        RECT 1389.290 57.745 1391.180 57.845 ;
        RECT 1389.290 56.160 1392.595 57.745 ;
        RECT 1389.310 56.145 1392.595 56.160 ;
        RECT 1389.310 53.110 1391.180 56.145 ;
        RECT 1202.430 0.195 1205.640 1.720 ;
        RECT 1202.430 0.120 1205.630 0.195 ;
      LAYER met5 ;
        RECT 1189.955 112.775 1193.395 112.900 ;
        RECT 1189.955 111.175 1510.590 112.775 ;
        RECT 1189.955 111.060 1193.395 111.175 ;
        RECT 1193.310 107.775 1196.750 107.800 ;
        RECT 1193.310 106.175 1510.590 107.775 ;
        RECT 1193.310 105.960 1196.750 106.175 ;
        RECT 1197.015 102.775 1200.455 102.915 ;
        RECT 1197.015 101.175 1510.590 102.775 ;
        RECT 1197.015 101.075 1200.455 101.175 ;
        RECT 1200.390 97.775 1203.830 97.840 ;
        RECT 1200.390 96.175 1510.590 97.775 ;
        RECT 1200.390 96.000 1203.830 96.175 ;
        RECT 1204.045 92.775 1207.485 92.860 ;
        RECT 1204.045 91.175 1510.590 92.775 ;
        RECT 1204.045 91.020 1207.485 91.175 ;
        RECT 1225.985 87.775 1229.425 87.830 ;
        RECT 1225.985 86.175 1510.590 87.775 ;
        RECT 1225.985 85.990 1229.425 86.175 ;
        RECT 1230.450 81.175 1510.590 82.775 ;
        RECT 1228.140 77.775 1231.580 77.860 ;
        RECT 1228.140 76.175 1510.590 77.775 ;
        RECT 1228.140 76.020 1231.580 76.175 ;
        RECT 1232.480 71.175 1510.590 72.775 ;
        RECT 1273.040 67.775 1276.480 67.825 ;
        RECT 1273.040 66.175 1510.590 67.775 ;
        RECT 1273.040 65.985 1276.480 66.175 ;
        RECT 1277.910 61.175 1510.590 62.775 ;
        RECT 1389.275 57.775 1392.715 57.865 ;
        RECT 1389.275 56.175 1510.590 57.775 ;
        RECT 1389.275 56.025 1392.715 56.175 ;
        RECT 1393.065 51.175 1510.590 52.775 ;
        RECT 1188.360 14.510 1191.800 15.680 ;
        RECT 0.000 13.840 1191.800 14.510 ;
        RECT 0.000 12.910 1190.170 13.840 ;
        RECT 1191.785 11.300 1195.225 12.175 ;
        RECT 0.000 10.335 1195.225 11.300 ;
        RECT 0.000 9.700 1193.700 10.335 ;
        RECT 1195.295 8.100 1198.735 8.730 ;
        RECT 0.000 6.890 1198.735 8.100 ;
        RECT 0.000 6.500 1197.020 6.890 ;
        RECT 1198.720 4.900 1202.160 5.285 ;
        RECT 0.000 3.445 1202.160 4.900 ;
        RECT 0.000 3.300 1201.100 3.445 ;
        RECT 1202.310 1.690 1205.750 1.840 ;
        RECT 0.000 0.090 1205.765 1.690 ;
        RECT 1202.310 0.000 1205.750 0.090 ;
  END
END analog_routes_bottom
END LIBRARY

