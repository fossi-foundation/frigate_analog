magic
tech sky130A
magscale 1 2
timestamp 1731205139
<< metal1 >>
rect 5574 19098 5682 19103
rect 5571 19077 5895 19098
rect 942 18822 1050 18823
rect 941 18804 1305 18822
rect 941 18525 961 18804
rect 1281 18525 1305 18804
rect 5571 18803 5586 19077
rect 5866 18803 5895 19077
rect 5571 18781 5895 18803
rect 10204 19081 10528 19103
rect 10204 18807 10219 19081
rect 10499 18807 10528 19081
rect 10204 18789 10528 18807
rect 14621 19082 14946 19103
rect 14621 18808 14646 19082
rect 14926 18808 14946 19082
rect 941 18505 1305 18525
rect -47 18373 251 18391
rect -47 18091 -27 18373
rect 228 18091 251 18373
rect -47 18072 251 18091
rect -47 4200 101 18072
rect 942 4226 1050 18505
rect 4584 18370 4908 18392
rect 4584 18096 4604 18370
rect 4884 18096 4908 18370
rect 4584 18075 4908 18096
rect 4585 4214 4733 18075
rect 5574 4192 5682 18781
rect 9214 18366 9538 18391
rect 9214 18092 9236 18366
rect 9516 18092 9538 18366
rect 9214 18074 9538 18092
rect 9217 4186 9365 18074
rect 10206 4250 10314 18789
rect 14621 18786 14946 18808
rect 13849 18367 14173 18388
rect 13849 18093 13867 18367
rect 14147 18093 14173 18367
rect 13849 18071 14173 18093
rect 13849 4204 13997 18071
rect 14838 4260 14946 18786
rect -288 -624 2270 -140
rect 2460 -624 6902 -140
rect 7092 -624 11534 -140
rect 11724 -624 16166 -140
rect 16356 -624 18156 -140
rect -288 -1326 3752 -842
rect 3920 -1326 8384 -842
rect 8552 -1326 13016 -842
rect 13184 -1326 17648 -842
rect 17816 -1326 18156 -842
<< via1 >>
rect 961 18525 1281 18804
rect 5586 18803 5866 19077
rect 10219 18807 10499 19081
rect 14646 18808 14926 19082
rect -27 18091 228 18373
rect 4604 18096 4884 18370
rect 9236 18092 9516 18366
rect 13867 18093 14147 18367
rect 2270 -624 2460 -140
rect 6902 -624 7092 -140
rect 11534 -624 11724 -140
rect 16166 -624 16356 -140
rect 3752 -1326 3920 -842
rect 8384 -1326 8552 -842
rect 13016 -1326 13184 -842
rect 17648 -1326 17816 -842
<< metal2 >>
rect 3112 19082 15058 19102
rect 3112 19081 14646 19082
rect 3112 19077 10219 19081
rect 3112 18822 5586 19077
rect -244 18804 5586 18822
rect -244 18525 961 18804
rect 1281 18803 5586 18804
rect 5866 18807 10219 19077
rect 10499 18808 14646 19081
rect 14926 18808 15058 19082
rect 10499 18807 15058 18808
rect 5866 18803 15058 18807
rect 1281 18784 15058 18803
rect 1281 18525 3520 18784
rect -244 18504 3520 18525
rect -244 18373 15058 18391
rect -244 18091 -27 18373
rect 228 18370 15058 18373
rect 228 18096 4604 18370
rect 4884 18367 15058 18370
rect 4884 18366 13867 18367
rect 4884 18096 9236 18366
rect 228 18092 9236 18096
rect 9516 18093 13867 18366
rect 14147 18093 15058 18367
rect 9516 18092 15058 18093
rect 228 18091 15058 18092
rect -244 18073 15058 18091
rect 6088 18012 6160 18026
rect 10714 18012 10778 18020
rect 4220 17976 6162 18012
rect 8852 17976 10794 18012
rect 13484 17976 15426 18012
rect 3168 17854 3600 17888
rect -412 17556 1425 17592
rect -412 -1454 -376 17556
rect -340 13464 1522 13500
rect -340 -1454 -304 13464
rect -268 8948 1538 8984
rect -268 -1454 -232 8948
rect -196 4432 1514 4468
rect -196 -1454 -160 4432
rect 2270 4233 2460 14643
rect 2608 13230 3040 14484
rect 3168 13030 3600 17320
rect 2608 8514 3040 9310
rect 3168 8482 3600 9976
rect 2608 3980 3040 4724
rect 3168 1376 3600 5456
rect 3752 4251 3920 14692
rect 2270 -140 2460 1168
rect 2270 -645 2460 -624
rect 3752 -842 3920 1146
rect 3752 -1338 3920 -1326
rect 4220 -1454 4256 17976
rect 6088 17762 6160 17976
rect 7800 17858 8232 17902
rect 8232 17404 8236 17556
rect 4292 13464 6154 13500
rect 4292 -1454 4328 13464
rect 4364 8948 6170 8984
rect 4364 -1454 4400 8948
rect 4436 4432 6146 4468
rect 4436 -1454 4472 4432
rect 6902 4227 7092 14615
rect 7240 14128 7672 14514
rect 7800 12994 8232 17324
rect 7800 8476 8232 9968
rect 7240 3990 7672 5202
rect 7800 3966 8232 5452
rect 8384 4238 8552 14648
rect 6902 -140 7092 1134
rect 6902 -645 7092 -624
rect 7800 -1436 8232 1356
rect 8384 -842 8552 1127
rect 8384 -1341 8552 -1326
rect 8852 -1454 8888 17976
rect 10714 17870 10778 17976
rect 12432 16949 12864 17218
rect 12864 16772 12868 16924
rect 12864 16456 12868 16608
rect 8924 13464 10786 13500
rect 8924 -1454 8960 13464
rect 8996 8948 10802 8984
rect 8996 -1454 9032 8948
rect 9068 4432 10778 4468
rect 9068 -1454 9104 4432
rect 11534 4227 11724 14623
rect 11874 13728 12304 14490
rect 12432 13030 12864 16415
rect 11872 8510 12304 9810
rect 12432 8516 12864 9980
rect 11872 3996 12304 4690
rect 12432 1410 12864 5454
rect 13016 4251 13184 14620
rect 11534 -140 11724 1109
rect 11534 -634 11724 -624
rect 13016 -842 13184 1105
rect 13484 462 13520 17976
rect 17064 16949 17496 17549
rect 13016 -1341 13184 -1326
rect 13244 426 13520 462
rect 13556 13464 15418 13500
rect 13244 -1454 13280 426
rect 13556 382 13592 13464
rect 13316 346 13592 382
rect 13628 8948 15434 8984
rect 13316 -1454 13352 346
rect 13628 308 13664 8948
rect 15350 8740 15434 8948
rect 13388 272 13664 308
rect 13700 4432 15410 4468
rect 13388 -1454 13424 272
rect 13700 226 13736 4432
rect 16166 4233 16356 14649
rect 16506 14128 16936 14478
rect 17064 12982 17496 16415
rect 16504 8506 16936 8794
rect 17064 8516 17496 9980
rect 16504 3982 16934 4688
rect 13460 190 13736 226
rect 13460 -1454 13496 190
rect 16166 -140 16356 1109
rect 16166 -634 16356 -624
rect 17064 -1404 17496 5464
rect 17648 4251 17816 14594
rect 17648 -842 17816 1105
rect 17648 -1341 17816 -1326
<< via2 >>
rect 3168 17320 3600 17854
rect 7800 17324 8232 17858
rect 12432 16415 12864 16949
rect 17064 16415 17496 16949
<< metal3 >>
rect 3126 17858 8298 17870
rect 3126 17854 7800 17858
rect 3126 17320 3168 17854
rect 3600 17324 7800 17854
rect 8232 17324 8298 17858
rect 3600 17320 8298 17324
rect 3126 17309 8298 17320
rect 12388 16949 17562 16962
rect 12388 16415 12432 16949
rect 12864 16415 17064 16949
rect 17496 16415 17562 16949
rect 12388 16401 17562 16415
rect -184 13749 19634 13877
rect -184 13237 19634 13365
rect -184 12725 19634 12853
rect -184 12213 19634 12341
rect -184 11701 19634 11829
rect -184 11189 19634 11317
rect -184 10677 19634 10805
rect -184 10165 19634 10293
rect -184 9653 19634 9781
rect -184 9141 19634 9269
rect -184 8629 19634 8757
rect -184 8117 19634 8245
rect -184 6581 19634 6709
rect -184 6069 19634 6197
rect -184 5557 19634 5685
rect -184 5045 19634 5173
<< metal4 >>
rect 7226 12286 7678 14176
rect 16510 12796 16934 14200
rect 2604 4610 3024 6146
rect 11878 4586 12306 6630
rect 16506 4598 16950 5608
use anablock_via_cut3  anablock_via_cut3_0
timestamp 1719104139
transform 0 1 9734 -1 0 10403
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_1
timestamp 1719104139
transform 0 1 -4162 -1 0 14918
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_2
timestamp 1719104139
transform 0 1 5102 -1 0 10403
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_3
timestamp 1719104139
transform 0 1 -4162 -1 0 10403
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_4
timestamp 1719104139
transform 0 1 -4162 -1 0 5888
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_5
timestamp 1719104139
transform 0 1 470 -1 0 5888
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_6
timestamp 1719104139
transform 0 1 5102 -1 0 5888
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_7
timestamp 1719104139
transform 0 1 9734 -1 0 5888
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_9
timestamp 1719104139
transform 0 1 9734 -1 0 14918
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_10
timestamp 1719104139
transform 0 1 5102 -1 0 14918
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_11
timestamp 1719104139
transform 0 1 470 -1 0 14918
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_12
timestamp 1719104139
transform 0 1 9734 -1 0 19433
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_13
timestamp 1719104139
transform 0 1 5102 -1 0 19433
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_14
timestamp 1719104139
transform 0 1 470 -1 0 19433
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_15
timestamp 1719104139
transform -1 0 2850 0 -1 23215
box 1426 5624 1624 5684
use anablock_via_cut3  anablock_via_cut3_16
timestamp 1719104139
transform 0 1 470 -1 0 10403
box 1426 5624 1624 5684
use cv3_via2_8cut  cv3_via2_8cut_0
timestamp 1719106786
transform 0 1 -45664 -1 0 11520
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_1
timestamp 1719106786
transform 0 1 -50298 -1 0 11536
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_2
timestamp 1719106786
transform 0 1 -45686 -1 0 15616
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_3
timestamp 1719106786
transform 0 1 -50312 -1 0 16648
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_4
timestamp 1719106786
transform 0 1 -45656 -1 0 17670
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_5
timestamp 1719106786
transform 0 1 -50298 -1 0 18686
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_7
timestamp 1719106786
transform 0 1 -50306 -1 0 20750
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_8
timestamp 1719106786
transform 0 1 -54920 -1 0 12044
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_9
timestamp 1719106786
transform 0 1 -59556 -1 0 11552
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_10
timestamp 1719106786
transform 0 1 -54928 -1 0 15116
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_11
timestamp 1719106786
transform 0 1 -59580 -1 0 16136
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_12
timestamp 1719106786
transform 0 1 -54926 -1 0 17168
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_13
timestamp 1719106786
transform 0 1 -59568 -1 0 18182
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_14
timestamp 1719106786
transform 0 1 -54942 -1 0 21142
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_15
timestamp 1719106786
transform 0 1 -59580 -1 0 20240
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_16
timestamp 1719106786
transform 0 1 -45674 -1 0 21142
box 6850 62208 6998 62544
use cv3_via3_10cut  cv3_via3_10cut_0
timestamp 1719433677
transform 1 0 -415714 0 1 -56350
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_1
timestamp 1719433677
transform 1 0 -429556 0 1 -65948
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_2
timestamp 1719433677
transform 1 0 -415726 0 1 -57774
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_3
timestamp 1719433677
transform 1 0 -424976 0 1 -56366
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_4
timestamp 1719433677
transform 1 0 -424992 0 1 -58290
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_5
timestamp 1719433677
transform 1 0 -429556 0 1 -64430
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_6
timestamp 1719433677
transform 1 0 -420330 0 1 -65948
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_7
timestamp 1719433677
transform 1 0 -420314 0 1 -63928
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_8
timestamp 1719433677
transform 1 0 -415680 0 1 -65958
box 431918 70502 432946 70630
use cv3_via3_10cut  cv3_via3_10cut_9
timestamp 1719433677
transform 1 0 -415690 0 1 -64948
box 431918 70502 432946 70630
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_1 ../dependencies/sky130_ef_ip__analog_switches/mag
array 0 3 -4515 0 3 -4632
timestamp 1731190834
transform 0 -1 3580 -1 0 4419
box -4 -600 3538 3648
<< labels >>
flabel metal3 18664 13813 18664 13813 0 FreeSans 960 0 0 0 right_instramp_p
flabel metal3 19082 13301 19082 13301 0 FreeSans 960 0 0 0 right_instramp_n
flabel metal3 19058 12785 19058 12785 0 FreeSans 960 0 0 0 right_lp_opamp_p
flabel metal3 18990 12271 18990 12271 0 FreeSans 960 0 0 0 right_lp_opamp_n
flabel metal3 18980 11767 18980 11767 0 FreeSans 960 0 0 0 right_hgbw_opamp_p
flabel metal3 19058 11249 19058 11249 0 FreeSans 960 0 0 0 right_hgbw_opamp_n
flabel metal3 19052 10741 19052 10741 0 FreeSans 960 0 0 0 left_hgbw_opamp_p
flabel metal3 19036 10235 19036 10235 0 FreeSans 960 0 0 0 left_hgbw_opamp_n
flabel metal3 19028 9715 19028 9715 0 FreeSans 960 0 0 0 left_lp_opamp_p
flabel metal3 18988 9213 18988 9213 0 FreeSans 960 0 0 0 left_lp_opamp_n
flabel metal3 19030 8695 19030 8695 0 FreeSans 960 0 0 0 left_instramp_p
flabel metal3 19014 8179 19014 8179 0 FreeSans 960 0 0 0 left_instramp_n
flabel metal3 18928 6649 18928 6649 0 FreeSans 960 0 0 0 ulpcomp_p
flabel metal3 18900 6131 18900 6131 0 FreeSans 960 0 0 0 ulpcomp_n
flabel metal3 18864 5619 18864 5619 0 FreeSans 960 0 0 0 comp_p
flabel metal3 18826 5107 18826 5107 0 FreeSans 960 0 0 0 comp_n
flabel metal2 17322 -1240 17322 -1240 0 FreeSans 1600 0 0 0 sio0
flabel metal1 223 -412 223 -412 0 FreeSans 1600 0 0 0 vdda0
flabel metal1 177 -1070 177 -1070 0 FreeSans 1600 0 0 0 vssa0
flabel metal2 8003 -1213 8003 -1213 0 FreeSans 1600 0 0 0 sio1
flabel metal2 2228 18211 2228 18211 0 FreeSans 1600 0 0 0 vssd0
flabel metal2 2284 18635 2284 18635 0 FreeSans 1600 0 0 0 vccd0
<< end >>
