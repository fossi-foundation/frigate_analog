magic
tech sky130A
magscale 1 2
timestamp 1717859832
<< metal3 >>
rect 30891 1250 31343 1272
rect 30891 1077 30920 1250
rect 31321 1077 31343 1250
rect 30891 1058 31343 1077
<< via3 >>
rect 30920 1077 31321 1250
<< metal4 >>
rect 571 2285 1571 2322
rect 571 2039 620 2285
rect 1539 2039 1571 2285
rect 571 285 1571 2039
rect 30223 1289 31376 1320
rect 30223 1029 30263 1289
rect 31001 1250 31376 1289
rect 31321 1077 31376 1250
rect 31001 1029 31376 1077
rect 30223 1000 31376 1029
rect 571 39 617 285
rect 1536 39 1571 285
rect 571 0 1571 39
<< via4 >>
rect 620 2039 1539 2285
rect 30263 1250 31001 1289
rect 30263 1077 30920 1250
rect 30920 1077 31001 1250
rect 30263 1029 31001 1077
rect 617 39 1536 285
<< metal5 >>
rect 0 2285 31032 2320
rect 0 2039 620 2285
rect 1539 2039 31032 2285
rect 0 2000 31032 2039
rect 298 1289 31038 1320
rect 298 1029 30263 1289
rect 31001 1029 31038 1289
rect 298 1000 31038 1029
rect 0 285 31032 320
rect 0 39 617 285
rect 1536 39 31032 285
rect 0 0 31032 39
<< properties >>
string FIXED_BBOX 0 0 31376 2322
string LEFclass COVER
<< end >>
