magic
tech sky130A
magscale 1 2
timestamp 1722440180
<< metal1 >>
rect 173599 41068 173605 41120
rect 173657 41111 173663 41120
rect 173657 41076 174299 41111
rect 173657 41068 173663 41076
rect 173946 38560 173952 38612
rect 174004 38604 174010 38612
rect 174004 38568 174350 38604
rect 174004 38560 174010 38568
rect 173946 17594 173952 17646
rect 174004 17638 174010 17646
rect 187560 17638 187596 18334
rect 174004 17602 187596 17638
rect 174004 17594 174010 17602
rect 173946 8514 173952 8522
rect 136762 8478 173952 8514
rect 173946 8470 173952 8478
rect 174004 8470 174010 8522
rect 170288 1969 179622 2005
rect 173600 1921 173606 1928
rect 170288 1885 173606 1921
rect 173600 1876 173606 1885
rect 173658 1876 173664 1928
<< via1 >>
rect 173605 41068 173657 41120
rect 173952 38560 174004 38612
rect 173952 17594 174004 17646
rect 173952 8470 174004 8522
rect 173606 1876 173658 1928
<< metal2 >>
rect 177261 50072 177461 50716
rect 177261 49872 180595 50072
rect 180395 47616 180595 49872
rect 173605 41120 173657 41126
rect 173605 41062 173657 41068
rect 150226 102 150262 8779
rect 150624 6969 150652 8744
rect 151033 7149 151061 8735
rect 151406 7299 151434 8758
rect 151795 7425 151823 8758
rect 152180 7580 152208 8726
rect 152550 8371 152578 8749
rect 152368 8343 152578 8371
rect 152180 7552 152284 7580
rect 151795 7397 152172 7425
rect 151406 7271 152060 7299
rect 151033 7121 151948 7149
rect 150624 6944 151836 6969
rect 150632 6941 151836 6944
rect 151808 0 151836 6941
rect 151920 0 151948 7121
rect 152032 0 152060 7271
rect 152144 0 152172 7397
rect 152256 0 152284 7552
rect 152368 0 152396 8343
rect 152930 8212 152958 8746
rect 152480 8184 152958 8212
rect 152480 0 152508 8184
rect 153314 8031 153342 8740
rect 152592 8003 153342 8031
rect 152592 0 152620 8003
rect 153692 7893 153720 8721
rect 152704 7865 153720 7893
rect 152704 0 152732 7865
rect 154055 7713 154083 8726
rect 152816 7685 154083 7713
rect 152816 0 152844 7685
rect 154451 7570 154479 8728
rect 152928 7542 154479 7570
rect 152928 0 152956 7542
rect 154817 7384 154845 8737
rect 153040 7356 154845 7384
rect 153040 0 153068 7356
rect 173614 1934 173649 41062
rect 173952 38612 174004 38618
rect 173952 38554 174004 38560
rect 173960 17652 173996 38554
rect 180312 35508 180512 36534
rect 179636 35408 180512 35508
rect 178943 31327 179043 32336
rect 179401 31323 179501 32963
rect 179636 31309 179736 35408
rect 173952 17646 174004 17652
rect 173952 17588 174004 17594
rect 173960 8528 173996 17588
rect 173952 8522 174004 8528
rect 173952 8464 174004 8470
rect 173606 1928 173658 1934
rect 173606 1870 173658 1876
rect 173614 1865 173649 1870
rect 179503 1794 179603 19922
rect 181186 19591 181682 20308
rect 182332 19596 182828 20072
rect 181176 19528 181713 19591
rect 181176 17927 181239 19528
rect 181638 17927 181713 19528
rect 181176 17835 181713 17927
rect 182326 19516 182863 19596
rect 182326 17915 182389 19516
rect 182788 17915 182863 19516
rect 182326 17840 182863 17915
<< via2 >>
rect 181239 17927 181638 19528
rect 182389 17915 182788 19516
<< metal3 >>
rect 174353 50716 174928 50826
rect 174354 47204 174432 50716
rect 174855 47204 174929 50716
rect 174354 47117 174929 47204
rect 170873 32879 179518 32941
rect 171672 32294 179056 32311
rect 171672 32194 171692 32294
rect 172672 32249 179056 32294
rect 172672 32194 172694 32249
rect 171672 32176 172694 32194
rect 181176 19528 181713 19591
rect 181176 17927 181239 19528
rect 181638 17927 181713 19528
rect 181176 17835 181713 17927
rect 182326 19516 182863 19596
rect 182326 17915 182389 19516
rect 182788 17915 182863 19516
rect 182326 17840 182863 17915
rect 136762 8396 190046 8406
rect 136762 8289 172516 8396
rect 172752 8289 190046 8396
rect 136762 8278 190046 8289
rect 136762 7932 190046 8132
rect 136762 7772 190046 7784
rect 136762 7665 172508 7772
rect 172744 7665 190046 7772
rect 136762 7656 190046 7665
rect 136762 7310 190046 7510
rect 136762 7151 190046 7162
rect 136762 7044 172508 7151
rect 172744 7044 190046 7151
rect 136762 7034 190046 7044
<< via3 >>
rect 153572 59658 155089 60010
rect 150103 59034 151655 59383
rect 174432 47204 174855 50716
rect 175531 36516 175764 38360
rect 171692 32194 172672 32294
rect 181239 17927 181638 19528
rect 182389 17915 182788 19516
rect 148574 9388 149640 9709
rect 155396 8804 156477 9135
rect 172516 8289 172752 8396
rect 172508 7665 172744 7772
rect 172508 7044 172744 7151
<< metal4 >>
rect 173626 69059 173943 69124
rect 173626 67913 173664 69059
rect 173901 67913 173943 69059
rect 153550 64947 155115 65290
rect 153550 63632 153658 64947
rect 155009 63632 155115 64947
rect 150076 62801 151681 63222
rect 150076 61486 150206 62801
rect 151557 61486 151681 62801
rect 150076 59383 151681 61486
rect 153550 60010 155115 63632
rect 153550 59658 153572 60010
rect 155089 59658 155115 60010
rect 153550 59623 155115 59658
rect 171674 62799 172694 63062
rect 171674 61472 171742 62799
rect 172605 61472 172694 62799
rect 150076 59034 150103 59383
rect 151655 59034 151681 59383
rect 150076 58995 151681 59034
rect 171674 32294 172694 61472
rect 173626 41840 173943 67913
rect 192853 69022 193914 69106
rect 192853 67944 192943 69022
rect 193812 67944 193914 69022
rect 175128 67097 175622 67169
rect 175128 65967 175168 67097
rect 175560 65967 175622 67097
rect 174354 64993 174929 65167
rect 174354 63571 174389 64993
rect 174887 63571 174929 64993
rect 174354 50716 174929 63571
rect 174354 47204 174432 50716
rect 174855 47204 174929 50716
rect 174354 47117 174929 47204
rect 175128 47028 175622 65967
rect 191197 64959 191960 65135
rect 191197 63620 191253 64959
rect 191878 63620 191960 64959
rect 188053 62857 188419 62965
rect 188053 61446 188099 62857
rect 188379 61446 188419 62857
rect 188053 47730 188419 61446
rect 173626 41523 175808 41840
rect 175491 38360 175808 41523
rect 175491 36516 175531 38360
rect 175764 36516 175808 38360
rect 175491 36484 175808 36516
rect 171674 32194 171692 32294
rect 172672 32194 172694 32294
rect 171674 25085 172694 32194
rect 191197 30792 191960 63620
rect 187453 30029 191960 30792
rect 171674 24065 175891 25085
rect 137668 8001 137905 9971
rect 138033 7312 138270 9992
rect 148524 9709 149674 9743
rect 148524 9388 148574 9709
rect 149640 9388 149674 9709
rect 148524 2174 149674 9388
rect 155339 9135 156521 9229
rect 155339 8804 155396 9135
rect 156477 8804 156521 9135
rect 155339 8769 156521 8804
rect 155356 4568 156515 8769
rect 166832 7336 167058 9972
rect 167200 7953 167426 9972
rect 172498 8396 172765 24065
rect 172498 8289 172516 8396
rect 172752 8289 172765 8396
rect 172498 7772 172765 8289
rect 172498 7665 172508 7772
rect 172744 7665 172765 7772
rect 172498 7151 172765 7665
rect 172498 7044 172508 7151
rect 172744 7044 172765 7151
rect 172498 7004 172765 7044
rect 181176 19528 181713 19591
rect 181176 17927 181239 19528
rect 181638 17927 181713 19528
rect 155356 3217 155461 4568
rect 156401 3217 156515 4568
rect 155356 3072 156515 3217
rect 181176 4639 181713 17927
rect 181176 3211 181249 4639
rect 181632 3211 181713 4639
rect 181176 3132 181713 3211
rect 182326 19516 182863 19596
rect 182326 17915 182389 19516
rect 182788 17915 182863 19516
rect 148524 823 148622 2174
rect 149562 823 149674 2174
rect 148524 580 149674 823
rect 182326 2221 182863 17915
rect 192853 4612 193914 67944
rect 192853 3207 192931 4612
rect 193816 3207 193914 4612
rect 192853 3072 193914 3207
rect 194710 67091 195771 67236
rect 194710 65970 194788 67091
rect 195667 65970 195771 67091
rect 182326 776 182365 2221
rect 182807 776 182863 2221
rect 182326 660 182863 776
rect 194710 2206 195771 65970
rect 194710 801 194793 2206
rect 195678 801 195771 2206
rect 194710 566 195771 801
<< via4 >>
rect 173664 67913 173901 69059
rect 153658 63632 155009 64947
rect 150206 61486 151557 62801
rect 171742 61472 172605 62799
rect 192943 67944 193812 69022
rect 175168 65967 175560 67097
rect 174389 63571 174887 64993
rect 191253 63620 191878 64959
rect 188099 61446 188379 62857
rect 155461 3217 156401 4568
rect 181249 3211 181632 4639
rect 148622 823 149562 2174
rect 192931 3207 193816 4612
rect 194788 65970 195667 67091
rect 182365 776 182807 2221
rect 194793 801 195678 2206
<< metal5 >>
rect 134778 69059 193994 69105
rect 134778 67913 173664 69059
rect 173901 69022 193994 69059
rect 173901 67944 192943 69022
rect 193812 67944 193994 69022
rect 173901 67913 193994 67944
rect 134778 67852 193994 67913
rect 134816 67097 195923 67168
rect 134816 65967 175168 67097
rect 175560 67091 195923 67097
rect 175560 65970 194788 67091
rect 195667 65970 195923 67091
rect 175560 65967 195923 65970
rect 134816 65915 195923 65967
rect 134593 64993 193084 65030
rect 134593 64947 174389 64993
rect 134593 63632 153658 64947
rect 155009 63632 174389 64947
rect 134593 63571 174389 63632
rect 174887 64959 193084 64993
rect 174887 63620 191253 64959
rect 191878 63620 193084 64959
rect 174887 63571 193084 63620
rect 134593 63536 193084 63571
rect 134806 62857 193297 62895
rect 134806 62801 188099 62857
rect 134806 61486 150206 62801
rect 151557 62799 188099 62801
rect 151557 61486 171742 62799
rect 134806 61472 171742 61486
rect 172605 61472 188099 62799
rect 134806 61446 188099 61472
rect 188379 61446 193297 62857
rect 134806 61401 193297 61446
rect 136826 4639 195936 4706
rect 136826 4568 181249 4639
rect 136826 3217 155461 4568
rect 156401 3217 181249 4568
rect 136826 3211 181249 3217
rect 181632 4612 195936 4639
rect 181632 3211 192931 4612
rect 136826 3207 192931 3211
rect 193816 3207 195936 4612
rect 136826 3138 195936 3207
rect 136826 2221 195980 2281
rect 136826 2174 182365 2221
rect 136826 823 148622 2174
rect 149562 823 182365 2174
rect 136826 776 182365 823
rect 182807 2206 195980 2221
rect 182807 801 194793 2206
rect 195678 801 195980 2206
rect 182807 776 195980 801
rect 136826 713 195980 776
use cv3_via2_8cut  cv3_via2_8cut_43
timestamp 1719106786
transform 1 0 172521 0 1 -29564
box 6850 62208 6998 62544
use cv3_via2_8cut  cv3_via2_8cut_44
timestamp 1719106786
transform 1 0 172065 0 1 -30221
box 6850 62208 6998 62544
use cv3_via3_30cut  cv3_via3_30cut_172
timestamp 1719173267
transform 1 0 -399491 0 1 -81257
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_173
timestamp 1719173267
transform 1 0 -399851 0 1 -81256
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_174
timestamp 1719173267
transform 1 0 -428657 0 1 -81255
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_175
timestamp 1719173267
transform 1 0 -429018 0 1 -81255
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_181
timestamp 1719173267
transform 0 1 45904 -1 0 574842
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_182
timestamp 1719173267
transform 0 1 76043 -1 0 574838
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_183
timestamp 1719173267
transform 0 1 75669 -1 0 574209
box 566656 91154 566956 91980
use cv3_via3_30cut  cv3_via3_30cut_184
timestamp 1719173267
transform 0 1 46273 -1 0 574213
box 566656 91154 566956 91980
use cv3_via_3cut  cv3_via_3cut_133
timestamp 1719452912
transform 1 0 168923 0 1 -105170
box 10601 106968 10663 107172
use sky130_ef_ip__ccomp3v_cl  sky130_ef_ip__ccomp3v_cl_1 ../ip/sky130_ef_ip__ccomp3v/mag
timestamp 1721179627
transform 0 1 177765 -1 0 31215
box -322 -2743 13304 10357
use sky130_ef_ip__cdac3v_12bit  sky130_ef_ip__cdac3v_12bit_0 ../ip/sky130_ef_ip__cdac3v_12bit/mag
timestamp 1722438219
transform 1 0 81345 0 -1 23288
box 52849 -36868 89580 14592
use sky130_ef_ip__samplehold  sky130_ef_ip__samplehold_0 ../ip/sky130_ef_ip__samplehold/mag
timestamp 1718244471
transform 1 0 173691 0 -1 48046
box 537 303 14883 11558
<< labels >>
flabel metal2 153040 0 153068 300 0 FreeSans 240 90 0 0 adc0_dac_val_11
port 640 nsew
flabel metal2 152928 0 152956 300 0 FreeSans 240 90 0 0 adc0_dac_val_10
port 641 nsew
flabel metal2 152816 0 152844 300 0 FreeSans 240 90 0 0 adc0_dac_val_9
port 642 nsew
flabel metal2 152704 0 152732 300 0 FreeSans 240 90 0 0 adc0_dac_val_8
port 643 nsew
flabel metal2 152592 0 152620 300 0 FreeSans 240 90 0 0 adc0_dac_val_7
port 644 nsew
flabel metal2 152480 0 152508 300 0 FreeSans 240 90 0 0 adc0_dac_val_6
port 645 nsew
flabel metal2 152368 0 152396 300 0 FreeSans 240 90 0 0 adc0_dac_val_5
port 646 nsew
flabel metal2 152256 0 152284 300 0 FreeSans 240 90 0 0 adc0_dac_val_4
port 647 nsew
flabel metal2 152144 0 152172 300 0 FreeSans 240 90 0 0 adc0_dac_val_3
port 648 nsew
flabel metal2 152032 0 152060 300 0 FreeSans 240 90 0 0 adc0_dac_val_2
port 649 nsew
flabel metal2 151920 0 151948 300 0 FreeSans 240 90 0 0 adc0_dac_val_1
port 650 nsew
flabel metal2 151808 0 151836 300 0 FreeSans 240 90 0 0 adc0_dac_val_0
port 651 nsew
flabel metal1 136762 8478 136866 8514 0 FreeSans 320 0 0 0 adc0_ena
port 652 nsew
flabel metal2 150226 102 150262 256 0 FreeSans 320 90 0 0 adc0_reset
port 653 nsew
flabel metal1 170288 1969 170425 2005 0 FreeSans 320 0 0 0 adc0_comp_out
port 654 nsew
flabel metal1 170288 1885 170426 1921 0 FreeSans 320 0 0 0 adc0_hold
port 656 nsew
flabel metal3 136762 7932 137018 8132 0 FreeSans 320 0 0 0 adc_vrefH
port 657 nsew
flabel metal3 136762 7310 137137 7510 0 FreeSans 320 0 0 0 adc_vrefL
port 658 nsew
flabel metal5 171792 3138 172938 4704 0 FreeSans 1600 0 0 0 vccd0
port 659 nsew
flabel metal5 171586 713 172629 2279 0 FreeSans 1600 0 0 0 vssd0
port 660 nsew
flabel metal3 174483 32902 174491 32911 0 FreeSans 800 0 0 0 adc_aval
flabel metal2 180040 35446 180040 35446 0 FreeSans 800 0 0 0 adc_sval
flabel metal2 177261 49872 177461 50716 0 FreeSans 800 90 0 0 adc0
port 662 nsew
flabel metal5 134965 61518 136829 62782 0 FreeSans 1600 0 0 0 vssa0
port 663 nsew
flabel metal5 134751 63658 136615 64922 0 FreeSans 1600 0 0 0 vdda0
port 664 nsew
<< end >>
