* NGSPICE file created from frigate_analog.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_g5v0d10v5_CPKWZQ w_n487_n797# a_29_n597# a_n287_n500# a_n229_n597#
+ a_229_n500# a_n29_n500#
X0 a_229_n500# a_29_n597# a_n29_n500# w_n487_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X1 a_n29_n500# a_n229_n597# a_n287_n500# w_n487_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_6THU7R a_n50_n597# a_50_n500# w_n308_n797# a_n108_n500#
X0 a_50_n500# a_n50_n597# a_n108_n500# w_n308_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_R6PXNO a_n287_n500# a_n487_n588# a_229_n500#
+ a_n545_n500# a_29_n588# a_n687_n722# a_n29_n500# a_487_n500# a_n229_n588# a_287_n588#
X0 a_487_n500# a_287_n588# a_229_n500# a_n687_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X1 a_229_n500# a_29_n588# a_n29_n500# a_n687_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_n29_n500# a_n229_n588# a_n287_n500# a_n687_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_n287_n500# a_n487_n588# a_n545_n500# a_n687_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_25MXQV a_n429_n588# a_29_n588# a_n487_n500# a_n629_n722#
+ a_n29_n500# a_429_n500#
X0 a_n29_n500# a_n429_n588# a_n487_n500# a_n629_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X1 a_429_n500# a_29_n588# a_n29_n500# a_n629_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_N7RQJ6 a_1261_n500# a_n1319_n500# a_1061_n588#
+ a_n287_n500# a_n1061_n500# a_n487_n588# a_745_n500# a_n1261_n588# a_545_n588# a_229_n500#
+ a_n545_n500# a_29_n588# a_1003_n500# a_n745_n588# a_n1461_n722# a_803_n588# a_n29_n500#
+ a_487_n500# a_n229_n588# a_n1003_n588# a_287_n588# a_n803_n500#
X0 a_n1061_n500# a_n1261_n588# a_n1319_n500# a_n1461_n722# sky130_fd_pr__nfet_05v0_nvt ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X1 a_1003_n500# a_803_n588# a_745_n500# a_n1461_n722# sky130_fd_pr__nfet_05v0_nvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_487_n500# a_287_n588# a_229_n500# a_n1461_n722# sky130_fd_pr__nfet_05v0_nvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_745_n500# a_545_n588# a_487_n500# a_n1461_n722# sky130_fd_pr__nfet_05v0_nvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a_1261_n500# a_1061_n588# a_1003_n500# a_n1461_n722# sky130_fd_pr__nfet_05v0_nvt ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X5 a_229_n500# a_29_n588# a_n29_n500# a_n1461_n722# sky130_fd_pr__nfet_05v0_nvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X6 a_n29_n500# a_n229_n588# a_n287_n500# a_n1461_n722# sky130_fd_pr__nfet_05v0_nvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X7 a_n545_n500# a_n745_n588# a_n803_n500# a_n1461_n722# sky130_fd_pr__nfet_05v0_nvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X8 a_n803_n500# a_n1003_n588# a_n1061_n500# a_n1461_n722# sky130_fd_pr__nfet_05v0_nvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X9 a_n287_n500# a_n487_n588# a_n545_n500# a_n1461_n722# sky130_fd_pr__nfet_05v0_nvt ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3P3PJP a_n50_n197# a_50_n100# w_n308_n397# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n308_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CBUN3Q a_29_n597# a_n287_n500# a_n229_n597# a_287_n597#
+ a_229_n500# w_n745_n797# a_n545_n500# a_n487_n597# a_n29_n500# a_487_n500#
X0 a_487_n500# a_287_n597# a_229_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X1 a_229_n500# a_29_n597# a_n29_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_n29_n500# a_n229_n597# a_n287_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_n287_n500# a_n487_n597# a_n545_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_5FCQ7L a_29_n597# a_n129_n597# a_129_n500# a_n29_n500#
+ w_n387_n797# a_n187_n500#
X0 a_129_n500# a_29_n597# a_n29_n500# w_n387_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X1 a_n29_n500# a_n129_n597# a_n187_n500# w_n387_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_VR3TSB a_50_n200# a_n242_n422# a_n108_n200# a_n50_n288#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n242_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_D5V3WB a_n429_n568# a_n487_n480# a_n29_n480#
+ a_29_n568# a_429_n480# a_n629_n702#
X0 a_429_n480# a_29_n568# a_n29_n480# a_n629_n702# sky130_fd_pr__nfet_g5v0d10v5 ad=1.392 pd=10.18 as=0.696 ps=5.09 w=4.8 l=2
X1 a_n29_n480# a_n429_n568# a_n487_n480# a_n629_n702# sky130_fd_pr__nfet_g5v0d10v5 ad=0.696 pd=5.09 as=1.392 ps=10.18 w=4.8 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TEGW2X a_n321_n472# a_29_n338# a_n29_n250# a_n129_n338#
+ a_n187_n250# a_129_n250#
X0 a_129_n250# a_29_n338# a_n29_n250# a_n321_n472# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=0.5
X1 a_n29_n250# a_n129_n338# a_n187_n250# a_n321_n472# sky130_fd_pr__nfet_g5v0d10v5 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=0.5
.ends

.subckt comparator_high_gain VDD VBN VSS VINP VOUT VINM DVDD ena3v3 w_355_n3243# DVSS
+ m2_4679_n3224#
XXM12 VDD m1_528_n2416# VDD m1_528_n2416# VDD m1_528_n2416# sky130_fd_pr__pfet_g5v0d10v5_CPKWZQ
XXM19 m1_4323_402# m1_3254_994# VDD VDD sky130_fd_pr__pfet_g5v0d10v5_6THU7R
XXM2 w_355_n3243# VINM w_355_n3243# m1_838_n2484# VINM w_355_n3243# m1_838_n2484#
+ m1_838_n2484# VINM VINM sky130_fd_pr__nfet_g5v0d10v5_R6PXNO
XXM3 VBN VBN w_355_n3243# VSS VSS w_355_n3243# sky130_fd_pr__nfet_g5v0d10v5_25MXQV
XXM5 m1_528_n2416# m1_528_n2416# VINM m1_528_n2416# m1_838_n2484# VINM m1_528_n2416#
+ VINM VINM m1_528_n2416# m1_838_n2484# VINM m1_838_n2484# VINM w_355_n3243# VINM
+ m1_838_n2484# m1_838_n2484# VINM VINM VINM m1_528_n2416# sky130_fd_pr__nfet_05v0_nvt_N7RQJ6
XXM8 ena3v3 VDD VDD m1_4323_402# sky130_fd_pr__pfet_g5v0d10v5_3P3PJP
XXM9 m1_528_n1044# m1_4323_402# m1_528_n1044# m1_528_n1044# m1_4323_402# VDD VDD m1_528_n1044#
+ VDD VDD sky130_fd_pr__pfet_g5v0d10v5_CBUN3Q
Xsky130_fd_pr__nfet_05v0_nvt_N7RQJ6_0 m1_528_n1044# m1_528_n1044# VINP m1_528_n1044#
+ m1_792_n1578# VINP m1_528_n1044# VINP VINP m1_528_n1044# m1_792_n1578# VINP m1_792_n1578#
+ VINP w_355_n3243# VINP m1_792_n1578# m1_792_n1578# VINP VINP VINP m1_528_n1044#
+ sky130_fd_pr__nfet_05v0_nvt_N7RQJ6
Xsky130_fd_pr__pfet_g5v0d10v5_5FCQ7L_0 m1_3254_994# m1_3254_994# VOUT DVDD VDD VOUT
+ sky130_fd_pr__pfet_g5v0d10v5_5FCQ7L
Xsky130_fd_pr__pfet_g5v0d10v5_CPKWZQ_0 VDD m1_528_n2416# VDD m1_528_n2416# VDD m1_528_n1044#
+ sky130_fd_pr__pfet_g5v0d10v5_CPKWZQ
XXM20 m1_3254_994# VSS VSS m1_4323_402# sky130_fd_pr__nfet_g5v0d10v5_VR3TSB
Xsky130_fd_pr__nfet_g5v0d10v5_R6PXNO_0 w_355_n3243# VINP w_355_n3243# m1_792_n1578#
+ VINP w_355_n3243# m1_792_n1578# m1_792_n1578# VINP VINP sky130_fd_pr__nfet_g5v0d10v5_R6PXNO
XXM10 VBN m1_4323_402# VSS VBN m1_4323_402# VSS sky130_fd_pr__nfet_g5v0d10v5_D5V3WB
XXM22 DVSS m1_3254_994# DVSS m1_3254_994# VOUT VOUT sky130_fd_pr__nfet_g5v0d10v5_TEGW2X
.ends

.subckt sky130_fd_pr__res_high_po_1p41_3L9D94 a_n141_2684# a_n897_2684# a_615_2684#
+ a_n141_n3116# a_n519_n3116# a_n1027_n3246# a_n897_n3116# a_237_n3116# a_615_n3116#
+ a_237_2684# a_n519_2684#
X0 a_n897_2684# a_n897_n3116# a_n1027_n3246# sky130_fd_pr__res_high_po_1p41 l=27
X1 a_615_2684# a_615_n3116# a_n1027_n3246# sky130_fd_pr__res_high_po_1p41 l=27
X2 a_n519_2684# a_n519_n3116# a_n1027_n3246# sky130_fd_pr__res_high_po_1p41 l=27
X3 a_n141_2684# a_n141_n3116# a_n1027_n3246# sky130_fd_pr__res_high_po_1p41 l=27
X4 a_237_2684# a_237_n3116# a_n1027_n3246# sky130_fd_pr__res_high_po_1p41 l=27
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_35MXHD a_n400_n722# a_200_n500# a_n258_n500#
+ a_n200_n588#
X0 a_200_n500# a_n200_n588# a_n258_n500# a_n400_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_VXYCT5 a_n200_n2097# a_200_n2000# w_n458_n2297#
+ a_n258_n2000#
X0 a_200_n2000# a_n200_n2097# a_n258_n2000# w_n458_n2297# sky130_fd_pr__pfet_g5v0d10v5 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_G59KN9 a_1500_n100# a_n1558_n100# w_n1758_n397#
+ a_n1500_n197#
X0 a_1500_n100# a_n1500_n197# a_n1558_n100# w_n1758_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=15
.ends

.subckt scomp_bias VDD VSS VBN ena3v3
XXR2 m1_3426_n1184# m1_4180_n1184# m1_785_3533# m1_3804_4616# m1_3804_4616# VSS VDD
+ m1_3048_4616# m1_3048_4616# m1_3426_n1184# m1_4180_n1184# sky130_fd_pr__res_high_po_1p41_3L9D94
XXM1 VSS m1_1110_n572# VSS VBN sky130_fd_pr__nfet_g5v0d10v5_35MXHD
XXM2 VSS VBN VSS VBN sky130_fd_pr__nfet_g5v0d10v5_35MXHD
XXM3 m1_785_3533# VDD VDD m1_1110_n572# sky130_fd_pr__pfet_g5v0d10v5_VXYCT5
XXM4 m1_1110_n572# m1_785_3533# VDD m1_1990_264# sky130_fd_pr__pfet_g5v0d10v5_VXYCT5
XXM5 VBN m1_785_3533# VDD VBN sky130_fd_pr__pfet_g5v0d10v5_G59KN9
XXM8 VSS m1_1990_264# VBN ena3v3 sky130_fd_pr__nfet_g5v0d10v5_35MXHD
.ends

.subckt sky130_fd_sc_hvl__lsbuflv2hv_1 A LVPWR VGND VPB VPWR X VPWR_uq0 VGND_uq0 VNB
X0 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2 X a_1711_885# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X3 X a_1711_885# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.12188 ps=1.075 w=0.75 l=0.5
X4 VGND_uq0 A a_404_1133# VNB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X5 a_1197_107# a_772_151# VGND_uq0 VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 VPWR_uq0 a_1197_107# a_504_1221# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X7 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X8 a_1197_107# a_772_151# VGND_uq0 VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X9 a_504_1221# a_404_1133# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X10 VGND a_404_1133# a_504_1221# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X11 a_772_151# a_404_1133# VGND_uq0 VNB sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X12 VGND_uq0 a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X13 LVPWR A a_404_1133# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X14 VPWR a_504_1221# a_1711_885# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X15 VGND a_504_1221# a_1711_885# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.12188 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X16 VGND_uq0 a_772_151# a_1197_107# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X17 a_772_151# a_404_1133# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X18 a_1197_107# a_772_151# VGND_uq0 VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X19 VPWR a_504_1221# a_1197_107# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1365 ps=1.49 w=0.42 l=1
.ends

.subckt sky130_fd_sc_hvl__diode_2 DIODE VGND VNB VPB VPWR
X0 VNB DIODE sky130_fd_pr__diode_pw2nd_11v0 perim=3.16e+06 area=6.072e+11
.ends

.subckt sky130_ef_ip__scomp3v VOUT VDD VINP VINM ENA DVDD w_6543_n2805# VSS w_7612_1960#
+ DVSS
Xx1 VDD x2/VBN VSS VINP VOUT VINM DVDD x3/X w_6543_n2805# DVSS VSS comparator_high_gain
Xx2 VDD VSS x2/VBN x3/X scomp_bias
Xx3 ENA DVDD DVSS VDD VDD x3/X VDD DVSS DVSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__diode_2_0 ENA DVSS DVSS VDD VDD sky130_fd_sc_hvl__diode_2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CVG6CD a_50_n400# w_n308_n697# a_n50_n464# a_n108_n400#
X0 a_50_n400# a_n50_n464# a_n108_n400# w_n308_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_W75H7K a_n4673_n1200# a_4873_n1200# a_2093_n1264#
+ a_n4099_n1264# w_n5131_n1497# a_4099_n1200# a_745_n1200# a_1577_n1264# a_803_n1264#
+ a_n745_n1264# a_n1003_n1264# a_n545_n1200# a_4157_n1264# a_n3583_n1264# a_3583_n1200#
+ a_1003_n1200# a_n3383_n1200# a_n2867_n1200# a_3641_n1264# a_n2293_n1264# a_2293_n1200#
+ a_n1577_n1200# a_n2093_n1200# a_n4931_n1200# a_2351_n1264# a_n1777_n1264# a_n4357_n1264#
+ a_1777_n1200# a_n29_n1200# a_n4157_n1200# a_1835_n1264# a_4357_n1200# a_n803_n1200#
+ a_4415_n1264# a_n3841_n1264# a_229_n1200# a_n3641_n1200# a_n229_n1264# a_3841_n1200#
+ a_1061_n1264# a_n3067_n1264# a_3067_n1200# a_3125_n1264# a_n2551_n1264# a_n2351_n1200#
+ a_2609_n1264# a_2551_n1200# a_n1835_n1200# a_n4615_n1264# a_4615_n1200# a_n4415_n1200#
+ a_1319_n1264# a_n1261_n1264# a_1261_n1200# a_n1061_n1200# a_3899_n1264# a_287_n1264#
+ a_n3325_n1264# a_n3125_n1200# a_n2809_n1264# a_3325_n1200# a_n2609_n1200# a_2809_n1200#
+ a_n2035_n1264# a_2035_n1200# a_n1519_n1264# a_1519_n1200# a_n1319_n1200# a_487_n1200#
+ a_n3899_n1200# a_4673_n1264# a_545_n1264# a_29_n1264# a_n487_n1264# a_n287_n1200#
+ a_3383_n1264# a_2867_n1264# a_n4873_n1264#
X0 a_1777_n1200# a_1577_n1264# a_1519_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X1 a_2809_n1200# a_2609_n1264# a_2551_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X2 a_n4157_n1200# a_n4357_n1264# a_n4415_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X3 a_1519_n1200# a_1319_n1264# a_1261_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X4 a_4873_n1200# a_4673_n1264# a_4615_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=1.74 ps=12.29 w=12 l=1
X5 a_3583_n1200# a_3383_n1264# a_3325_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X6 a_4615_n1200# a_4415_n1264# a_4357_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X7 a_n2867_n1200# a_n3067_n1264# a_n3125_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X8 a_487_n1200# a_287_n1264# a_229_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X9 a_2293_n1200# a_2093_n1264# a_2035_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X10 a_3325_n1200# a_3125_n1264# a_3067_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X11 a_n287_n1200# a_n487_n1264# a_n545_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X12 a_n2609_n1200# a_n2809_n1264# a_n2867_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X13 a_n1577_n1200# a_n1777_n1264# a_n1835_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X14 a_n29_n1200# a_n229_n1264# a_n287_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X15 a_n4673_n1200# a_n4873_n1264# a_n4931_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=3.48 ps=24.58 w=12 l=1
X16 a_2035_n1200# a_1835_n1264# a_1777_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X17 a_n1319_n1200# a_n1519_n1264# a_n1577_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X18 a_n4415_n1200# a_n4615_n1264# a_n4673_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X19 a_n3383_n1200# a_n3583_n1264# a_n3641_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X20 a_n3125_n1200# a_n3325_n1264# a_n3383_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X21 a_3841_n1200# a_3641_n1264# a_3583_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X22 a_n2093_n1200# a_n2293_n1264# a_n2351_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X23 a_745_n1200# a_545_n1264# a_487_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X24 a_n1835_n1200# a_n2035_n1264# a_n2093_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X25 a_2551_n1200# a_2351_n1264# a_2293_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X26 a_1261_n1200# a_1061_n1264# a_1003_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X27 a_n545_n1200# a_n745_n1264# a_n803_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X28 a_229_n1200# a_29_n1264# a_n29_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X29 a_4099_n1200# a_3899_n1264# a_3841_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X30 a_n3641_n1200# a_n3841_n1264# a_n3899_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X31 a_n2351_n1200# a_n2551_n1264# a_n2609_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X32 a_1003_n1200# a_803_n1264# a_745_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X33 a_n3899_n1200# a_n4099_n1264# a_n4157_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X34 a_n1061_n1200# a_n1261_n1264# a_n1319_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X35 a_4357_n1200# a_4157_n1264# a_4099_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X36 a_n803_n1200# a_n1003_n1264# a_n1061_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X37 a_3067_n1200# a_2867_n1264# a_2809_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_WKXP7K a_n4673_n1200# a_4873_n1200# a_4931_n1264#
+ a_2093_n1264# a_n4099_n1264# a_4099_n1200# a_745_n1200# a_1577_n1264# a_803_n1264#
+ a_n745_n1264# a_n1003_n1264# a_n545_n1200# a_4157_n1264# a_n3583_n1264# a_3583_n1200#
+ a_1003_n1200# a_n3383_n1200# a_n2867_n1200# a_3641_n1264# a_n2293_n1264# a_2293_n1200#
+ a_n1577_n1200# a_n2093_n1200# a_n4931_n1200# a_2351_n1264# a_n1777_n1264# a_n4357_n1264#
+ a_1777_n1200# a_n29_n1200# a_n4157_n1200# a_1835_n1264# a_4357_n1200# a_n803_n1200#
+ a_4415_n1264# a_n3841_n1264# a_229_n1200# a_n3641_n1200# a_n229_n1264# a_3841_n1200#
+ a_1061_n1264# a_n3067_n1264# a_3067_n1200# a_3125_n1264# a_n2551_n1264# a_n2351_n1200#
+ a_2609_n1264# a_n5131_n1264# w_n5389_n1497# a_5131_n1200# a_2551_n1200# a_n1835_n1200#
+ a_n4615_n1264# a_4615_n1200# a_n4415_n1200# a_1319_n1264# a_n1261_n1264# a_1261_n1200#
+ a_n1061_n1200# a_3899_n1264# a_287_n1264# a_n3325_n1264# a_n3125_n1200# a_n2809_n1264#
+ a_3325_n1200# a_n2609_n1200# a_2809_n1200# a_n2035_n1264# a_2035_n1200# a_n1519_n1264#
+ a_1519_n1200# a_n1319_n1200# a_487_n1200# a_n3899_n1200# a_4673_n1264# a_545_n1264#
+ a_29_n1264# a_n487_n1264# a_n287_n1200# a_3383_n1264# a_n5189_n1200# a_2867_n1264#
+ a_n4873_n1264#
X0 a_1777_n1200# a_1577_n1264# a_1519_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X1 a_2809_n1200# a_2609_n1264# a_2551_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X2 a_n4157_n1200# a_n4357_n1264# a_n4415_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X3 a_1519_n1200# a_1319_n1264# a_1261_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X4 a_4873_n1200# a_4673_n1264# a_4615_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X5 a_3583_n1200# a_3383_n1264# a_3325_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X6 a_4615_n1200# a_4415_n1264# a_4357_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X7 a_n2867_n1200# a_n3067_n1264# a_n3125_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X8 a_487_n1200# a_287_n1264# a_229_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X9 a_2293_n1200# a_2093_n1264# a_2035_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X10 a_3325_n1200# a_3125_n1264# a_3067_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X11 a_n287_n1200# a_n487_n1264# a_n545_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X12 a_n2609_n1200# a_n2809_n1264# a_n2867_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X13 a_n1577_n1200# a_n1777_n1264# a_n1835_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X14 a_n29_n1200# a_n229_n1264# a_n287_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X15 a_n4673_n1200# a_n4873_n1264# a_n4931_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X16 a_2035_n1200# a_1835_n1264# a_1777_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X17 a_n1319_n1200# a_n1519_n1264# a_n1577_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X18 a_5131_n1200# a_4931_n1264# a_4873_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=1.74 ps=12.29 w=12 l=1
X19 a_n4415_n1200# a_n4615_n1264# a_n4673_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X20 a_n3383_n1200# a_n3583_n1264# a_n3641_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X21 a_n3125_n1200# a_n3325_n1264# a_n3383_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X22 a_3841_n1200# a_3641_n1264# a_3583_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X23 a_n2093_n1200# a_n2293_n1264# a_n2351_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X24 a_745_n1200# a_545_n1264# a_487_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X25 a_n1835_n1200# a_n2035_n1264# a_n2093_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X26 a_2551_n1200# a_2351_n1264# a_2293_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X27 a_n4931_n1200# a_n5131_n1264# a_n5189_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=3.48 ps=24.58 w=12 l=1
X28 a_1261_n1200# a_1061_n1264# a_1003_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X29 a_n545_n1200# a_n745_n1264# a_n803_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X30 a_229_n1200# a_29_n1264# a_n29_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X31 a_4099_n1200# a_3899_n1264# a_3841_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X32 a_n3641_n1200# a_n3841_n1264# a_n3899_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X33 a_n2351_n1200# a_n2551_n1264# a_n2609_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X34 a_1003_n1200# a_803_n1264# a_745_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X35 a_n3899_n1200# a_n4099_n1264# a_n4157_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X36 a_n1061_n1200# a_n1261_n1264# a_n1319_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X37 a_4357_n1200# a_4157_n1264# a_4099_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X38 a_n803_n1200# a_n1003_n1264# a_n1061_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X39 a_3067_n1200# a_2867_n1264# a_2809_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_AALY9X c1_n5378_n3920# c1_5116_n3920# m3_8574_n3960#
+ c1_n1880_n3920# c1_1618_n3920# m3_n5418_n3960# m3_n1920_n3960# m3_5076_n3960# c1_n8876_n3920#
+ c1_8614_n3920# m3_1578_n3960# m3_n8916_n3960#
X0 c1_5116_n3920# m3_5076_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X1 c1_1618_n3920# m3_1578_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X2 c1_8614_n3920# m3_8574_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X3 c1_n5378_n3920# m3_n5418_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X4 c1_n8876_n3920# m3_n8916_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X5 c1_n5378_n3920# m3_n5418_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X6 c1_n1880_n3920# m3_n1920_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X7 c1_1618_n3920# m3_1578_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X8 c1_n8876_n3920# m3_n8916_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X9 c1_n5378_n3920# m3_n5418_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X10 c1_n8876_n3920# m3_n8916_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X11 c1_1618_n3920# m3_1578_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X12 c1_8614_n3920# m3_8574_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X13 c1_5116_n3920# m3_5076_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X14 c1_5116_n3920# m3_5076_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X15 c1_8614_n3920# m3_8574_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X16 c1_n1880_n3920# m3_n1920_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X17 c1_n1880_n3920# m3_n1920_n3960# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
.ends

.subckt sky130_fd_pr__nfet_01v8_6H2JYD a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CTEUHA a_50_n200# a_n242_n422# a_n108_n200# a_n50_n288#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n242_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_HQ4STX w_n358_n597# a_n158_n300# a_n100_n364#
+ a_100_n300#
X0 a_100_n300# a_n100_n364# a_n158_n300# w_n358_n597# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UKVZ7J a_1519_n450# a_n803_n450# a_n2093_n450#
+ a_n2551_n505# a_1261_n450# a_29_n505# a_n1777_n505# a_n3067_n505# a_n1319_n450#
+ a_n287_n450# a_n1061_n450# a_2867_n505# a_n745_n505# a_2809_n450# a_803_n505# a_n2035_n505#
+ a_745_n450# a_n3383_n450# a_2551_n450# a_3125_n505# a_1835_n505# a_3067_n450# a_1777_n450#
+ a_n2609_n450# a_n229_n505# a_n1003_n505# a_n2351_n450# a_287_n505# a_2093_n505#
+ a_229_n450# a_n1577_n450# a_n3325_n505# a_2035_n450# a_1319_n505# a_n545_n450# a_1061_n505#
+ a_n2293_n505# a_n3517_n672# a_1003_n450# a_n1519_n505# a_n2867_n450# a_n487_n505#
+ a_3325_n450# a_n1261_n505# a_2609_n505# a_n29_n450# a_545_n505# a_487_n450# a_2351_n505#
+ a_2293_n450# a_n1835_n450# a_n3125_n450# a_1577_n505# a_n2809_n505#
X0 a_n2093_n450# a_n2293_n505# a_n2351_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X1 a_229_n450# a_29_n505# a_n29_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X2 a_n29_n450# a_n229_n505# a_n287_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X3 a_3067_n450# a_2867_n505# a_2809_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X4 a_n1319_n450# a_n1519_n505# a_n1577_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X5 a_2551_n450# a_2351_n505# a_2293_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X6 a_n3125_n450# a_n3325_n505# a_n3383_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=1
X7 a_n545_n450# a_n745_n505# a_n803_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X8 a_n287_n450# a_n487_n505# a_n545_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X9 a_2293_n450# a_2093_n505# a_2035_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X10 a_n2867_n450# a_n3067_n505# a_n3125_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X11 a_n803_n450# a_n1003_n505# a_n1061_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X12 a_n1577_n450# a_n1777_n505# a_n1835_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X13 a_1519_n450# a_1319_n505# a_1261_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X14 a_n1061_n450# a_n1261_n505# a_n1319_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X15 a_3325_n450# a_3125_n505# a_3067_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=1
X16 a_1003_n450# a_803_n505# a_745_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X17 a_745_n450# a_545_n505# a_487_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X18 a_487_n450# a_287_n505# a_229_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X19 a_1777_n450# a_1577_n505# a_1519_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X20 a_2035_n450# a_1835_n505# a_1777_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X21 a_n2609_n450# a_n2809_n505# a_n2867_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X22 a_1261_n450# a_1061_n505# a_1003_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X23 a_n1835_n450# a_n2035_n505# a_n2093_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X24 a_2809_n450# a_2609_n505# a_2551_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X25 a_n2351_n450# a_n2551_n505# a_n2609_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_USXRNR a_1448_n255# a_1190_n255# a_358_n200#
+ a_n1648_n255# a_n1706_n200# a_100_n200# a_n674_n200# a_n616_n255# a_n1390_n255#
+ a_674_n255# a_1132_n200# a_n158_n200# a_158_n255# a_616_n200# a_n874_n255# a_n932_n200#
+ a_1648_n200# a_932_n255# a_1390_n200# a_n1448_n200# a_n358_n255# a_n416_n200# a_n1190_n200#
+ a_n1132_n255# a_874_n200# a_416_n255# a_n100_n255# a_n1840_n422#
X0 a_874_n200# a_674_n255# a_616_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_1132_n200# a_932_n255# a_874_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_1390_n200# a_1190_n255# a_1132_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_100_n200# a_n100_n255# a_n158_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_n416_n200# a_n616_n255# a_n674_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_n158_n200# a_n358_n255# a_n416_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_n1448_n200# a_n1648_n255# a_n1706_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X7 a_n1190_n200# a_n1390_n255# a_n1448_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_n674_n200# a_n874_n255# a_n932_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_n932_n200# a_n1132_n255# a_n1190_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_358_n200# a_158_n255# a_100_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_616_n200# a_416_n255# a_358_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X12 a_1648_n200# a_1448_n255# a_1390_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AUMBFF a_n2035_n2564# a_n1519_n2564# a_2035_n2500#
+ a_n1319_n2500# a_1519_n2500# a_n3899_n2500# a_487_n2500# a_545_n2564# a_29_n2564#
+ a_n487_n2564# a_n287_n2500# a_3383_n2564# a_2867_n2564# a_2093_n2564# a_n4099_n2564#
+ a_745_n2500# a_1577_n2564# a_803_n2564# a_n1003_n2564# w_n4615_n2797# a_4099_n2500#
+ a_n545_n2500# a_4157_n2564# a_n745_n2564# a_n3583_n2564# a_1003_n2500# a_n3383_n2500#
+ a_3583_n2500# a_n2867_n2500# a_3641_n2564# a_n2293_n2564# a_2293_n2500# a_n2093_n2500#
+ a_n1777_n2564# a_1777_n2500# a_n29_n2500# a_n1577_n2500# a_n4157_n2500# a_2351_n2564#
+ a_n4357_n2564# a_4357_n2500# a_1835_n2564# a_229_n2500# a_n803_n2500# a_n229_n2564#
+ a_n3841_n2564# a_3841_n2500# a_n3641_n2500# a_1061_n2564# a_n3067_n2564# a_3067_n2500#
+ a_3125_n2564# a_n2551_n2564# a_n2351_n2500# a_2609_n2564# a_2551_n2500# a_n1835_n2500#
+ a_n4415_n2500# a_1319_n2564# a_n1261_n2564# a_1261_n2500# a_n1061_n2500# a_3899_n2564#
+ a_n3125_n2500# a_287_n2564# a_n2809_n2564# a_n3325_n2564# a_3325_n2500# a_n2609_n2500#
+ a_2809_n2500#
X0 a_3067_n2500# a_2867_n2564# a_2809_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X1 a_2809_n2500# a_2609_n2564# a_2551_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X2 a_1777_n2500# a_1577_n2564# a_1519_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X3 a_1519_n2500# a_1319_n2564# a_1261_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X4 a_n4157_n2500# a_n4357_n2564# a_n4415_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=7.25 ps=50.58 w=25 l=1
X5 a_n2867_n2500# a_n3067_n2564# a_n3125_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X6 a_3583_n2500# a_3383_n2564# a_3325_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X7 a_487_n2500# a_287_n2564# a_229_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X8 a_2293_n2500# a_2093_n2564# a_2035_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X9 a_3325_n2500# a_3125_n2564# a_3067_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X10 a_n287_n2500# a_n487_n2564# a_n545_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X11 a_n2609_n2500# a_n2809_n2564# a_n2867_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X12 a_n1577_n2500# a_n1777_n2564# a_n1835_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X13 a_n29_n2500# a_n229_n2564# a_n287_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X14 a_2035_n2500# a_1835_n2564# a_1777_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X15 a_n1319_n2500# a_n1519_n2564# a_n1577_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X16 a_n3383_n2500# a_n3583_n2564# a_n3641_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X17 a_3841_n2500# a_3641_n2564# a_3583_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X18 a_n3125_n2500# a_n3325_n2564# a_n3383_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X19 a_n2093_n2500# a_n2293_n2564# a_n2351_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X20 a_745_n2500# a_545_n2564# a_487_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X21 a_n1835_n2500# a_n2035_n2564# a_n2093_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X22 a_2551_n2500# a_2351_n2564# a_2293_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X23 a_1261_n2500# a_1061_n2564# a_1003_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X24 a_n545_n2500# a_n745_n2564# a_n803_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X25 a_229_n2500# a_29_n2564# a_n29_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X26 a_4099_n2500# a_3899_n2564# a_3841_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X27 a_n3641_n2500# a_n3841_n2564# a_n3899_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X28 a_n2351_n2500# a_n2551_n2564# a_n2609_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X29 a_1003_n2500# a_803_n2564# a_745_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X30 a_n3899_n2500# a_n4099_n2564# a_n4157_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X31 a_n1061_n2500# a_n1261_n2564# a_n1319_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X32 a_4357_n2500# a_4157_n2564# a_4099_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=7.25 pd=50.58 as=3.625 ps=25.29 w=25 l=1
X33 a_n803_n2500# a_n1003_n2564# a_n1061_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_25PWK4 a_n148_n148# a_n46_n46#
X0 a_n148_n148# a_n46_n46# sky130_fd_pr__diode_pw2nd_05v5 perim=1.84e+06 area=2.116e+11
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QL2RRT a_29_n664# a_n1777_n664# a_n2351_n600#
+ a_n745_n664# a_229_n600# a_n1577_n600# a_2867_n664# a_2035_n600# a_803_n664# a_n2035_n664#
+ a_n545_n600# a_3125_n664# a_1835_n664# a_1003_n600# a_n229_n664# w_n3583_n897# a_287_n664#
+ a_n1003_n664# a_n2867_n600# a_3325_n600# a_2093_n664# a_n3325_n664# a_n29_n600#
+ a_487_n600# a_1319_n664# a_2293_n600# a_n3125_n600# a_n2293_n664# a_n1835_n600#
+ a_1061_n664# a_n803_n600# a_1519_n600# a_n2093_n600# a_n1519_n664# a_1261_n600#
+ a_n487_n664# a_n1261_n664# a_2609_n664# a_545_n664# a_n1319_n600# a_n287_n600# a_n1061_n600#
+ a_2351_n664# a_2809_n600# a_1577_n664# a_745_n600# a_n3383_n600# a_n2809_n664# a_2551_n600#
+ a_n2551_n664# a_3067_n600# a_1777_n600# a_n2609_n600# a_n3067_n664#
X0 a_2809_n600# a_2609_n664# a_2551_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X1 a_n2351_n600# a_n2551_n664# a_n2609_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X2 a_n2093_n600# a_n2293_n664# a_n2351_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X3 a_229_n600# a_29_n664# a_n29_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X4 a_n29_n600# a_n229_n664# a_n287_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X5 a_3067_n600# a_2867_n664# a_2809_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X6 a_n1319_n600# a_n1519_n664# a_n1577_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X7 a_2551_n600# a_2351_n664# a_2293_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X8 a_n3125_n600# a_n3325_n664# a_n3383_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=1
X9 a_n545_n600# a_n745_n664# a_n803_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X10 a_n287_n600# a_n487_n664# a_n545_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X11 a_2293_n600# a_2093_n664# a_2035_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X12 a_n2867_n600# a_n3067_n664# a_n3125_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X13 a_n803_n600# a_n1003_n664# a_n1061_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X14 a_n1577_n600# a_n1777_n664# a_n1835_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X15 a_1519_n600# a_1319_n664# a_1261_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X16 a_n1061_n600# a_n1261_n664# a_n1319_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X17 a_3325_n600# a_3125_n664# a_3067_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=1
X18 a_1003_n600# a_803_n664# a_745_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X19 a_745_n600# a_545_n664# a_487_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X20 a_487_n600# a_287_n664# a_229_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X21 a_2035_n600# a_1835_n664# a_1777_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X22 a_n2609_n600# a_n2809_n664# a_n2867_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X23 a_1777_n600# a_1577_n664# a_1519_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X24 a_1261_n600# a_1061_n664# a_1003_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X25 a_n1835_n600# a_n2035_n664# a_n2093_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_AALY9W c2_3778_n4000# c2_280_n4000# m4_n6796_n4080#
+ m4_7196_n4080# c2_n6716_n4000# m4_n10294_n4080# m4_3698_n4080# m4_n3298_n4080# c2_n10214_n4000#
+ m4_200_n4080# c2_7276_n4000# c2_n3218_n4000#
X0 c2_7276_n4000# m4_7196_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X1 c2_280_n4000# m4_200_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X2 c2_n3218_n4000# m4_n3298_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X3 c2_280_n4000# m4_200_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X4 c2_n6716_n4000# m4_n6796_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X5 c2_3778_n4000# m4_3698_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X6 c2_280_n4000# m4_200_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X7 c2_3778_n4000# m4_3698_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X8 c2_n10214_n4000# m4_n10294_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X9 c2_n10214_n4000# m4_n10294_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X10 c2_7276_n4000# m4_7196_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X11 c2_n6716_n4000# m4_n6796_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X12 c2_3778_n4000# m4_3698_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X13 c2_n3218_n4000# m4_n3298_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X14 c2_n10214_n4000# m4_n10294_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X15 c2_n6716_n4000# m4_n6796_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X16 c2_n3218_n4000# m4_n3298_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
X17 c2_7276_n4000# m4_7196_n4080# sky130_fd_pr__cap_mim_m3_2 l=12 w=12
.ends

.subckt sky130_fd_pr__pfet_01v8_U4BBJH a_15_n200# w_n211_n419# a_n33_n297# a_n73_n200#
X0 a_15_n200# a_n33_n297# a_n73_n200# w_n211_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_B3XH3Z a_1519_n450# a_n803_n450# a_n2093_n450#
+ a_n2551_n505# a_1261_n450# a_29_n505# a_n1777_n505# a_n3067_n505# a_n1319_n450#
+ a_3641_n505# a_3583_n450# a_n4033_n672# a_n287_n450# a_n1061_n450# a_2867_n505#
+ a_n745_n505# a_2809_n450# a_803_n505# a_n2035_n505# a_745_n450# a_n3383_n450# a_n3841_n505#
+ a_2551_n450# a_3125_n505# a_1835_n505# a_3067_n450# a_1777_n450# a_n2609_n450# a_n229_n505#
+ a_n1003_n505# a_n2351_n450# a_287_n505# a_2093_n505# a_229_n450# a_n1577_n450# a_n3325_n505#
+ a_2035_n450# a_3841_n450# a_1319_n505# a_n545_n450# a_n3899_n450# a_1061_n505# a_n2293_n505#
+ a_1003_n450# a_n3641_n450# a_3383_n505# a_n1519_n505# a_n2867_n450# a_n487_n505#
+ a_3325_n450# a_n1261_n505# a_2609_n505# a_n29_n450# a_545_n505# a_487_n450# a_2351_n505#
+ a_n3583_n505# a_2293_n450# a_n1835_n450# a_n3125_n450# a_1577_n505# a_n2809_n505#
X0 a_n2093_n450# a_n2293_n505# a_n2351_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X1 a_229_n450# a_29_n505# a_n29_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X2 a_n29_n450# a_n229_n505# a_n287_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X3 a_3067_n450# a_2867_n505# a_2809_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X4 a_n1319_n450# a_n1519_n505# a_n1577_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X5 a_2551_n450# a_2351_n505# a_2293_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X6 a_n3125_n450# a_n3325_n505# a_n3383_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X7 a_n545_n450# a_n745_n505# a_n803_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X8 a_n287_n450# a_n487_n505# a_n545_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X9 a_2293_n450# a_2093_n505# a_2035_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X10 a_n2867_n450# a_n3067_n505# a_n3125_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X11 a_n803_n450# a_n1003_n505# a_n1061_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X12 a_n3641_n450# a_n3841_n505# a_n3899_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=1
X13 a_n3383_n450# a_n3583_n505# a_n3641_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X14 a_n1577_n450# a_n1777_n505# a_n1835_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X15 a_1519_n450# a_1319_n505# a_1261_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X16 a_n1061_n450# a_n1261_n505# a_n1319_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X17 a_3325_n450# a_3125_n505# a_3067_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X18 a_1003_n450# a_803_n505# a_745_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X19 a_745_n450# a_545_n505# a_487_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X20 a_487_n450# a_287_n505# a_229_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X21 a_1777_n450# a_1577_n505# a_1519_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X22 a_2035_n450# a_1835_n505# a_1777_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X23 a_3841_n450# a_3641_n505# a_3583_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=1
X24 a_n2609_n450# a_n2809_n505# a_n2867_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X25 a_3583_n450# a_3383_n505# a_3325_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X26 a_1261_n450# a_1061_n505# a_1003_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X27 a_n1835_n450# a_n2035_n505# a_n2093_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X28 a_2809_n450# a_2609_n505# a_2551_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X29 a_n2351_n450# a_n2551_n505# a_n2609_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QTY6KC a_287_n464# a_n1003_n464# a_487_n400#
+ a_n29_n400# a_1319_n464# w_n1777_n697# a_1061_n464# a_1519_n400# a_n803_n400# a_n1519_n464#
+ a_1261_n400# a_n487_n464# a_n1261_n464# a_n1319_n400# a_545_n464# a_n287_n400# a_n1061_n400#
+ a_745_n400# a_29_n464# a_n745_n464# a_229_n400# a_n1577_n400# a_803_n464# a_n545_n400#
+ a_1003_n400# a_n229_n464#
X0 a_n1319_n400# a_n1519_n464# a_n1577_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X1 a_n545_n400# a_n745_n464# a_n803_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X2 a_n803_n400# a_n1003_n464# a_n1061_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 a_n287_n400# a_n487_n464# a_n545_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X4 a_1519_n400# a_1319_n464# a_1261_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X5 a_n1061_n400# a_n1261_n464# a_n1319_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X6 a_1003_n400# a_803_n464# a_745_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X7 a_487_n400# a_287_n464# a_229_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X8 a_745_n400# a_545_n464# a_487_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X9 a_1261_n400# a_1061_n464# a_1003_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X10 a_229_n400# a_29_n464# a_n29_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X11 a_n29_n400# a_n229_n464# a_n287_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_2B7385 a_1261_n800# a_n1319_n800# a_1835_n855#
+ a_n287_n800# a_n229_n855# a_n1061_n800# a_287_n855# a_n1003_n855# a_2093_n855# a_745_n800#
+ a_1319_n855# a_1777_n800# a_n2293_n855# a_n2351_n800# a_1061_n855# a_229_n800# a_2035_n800#
+ a_n1577_n800# a_n1519_n855# a_n487_n855# a_n1261_n855# a_n545_n800# a_545_n855#
+ a_1003_n800# a_1577_n855# a_n2485_n1022# a_n29_n800# a_487_n800# a_2293_n800# a_29_n855#
+ a_n1777_n855# a_n1835_n800# a_n745_n855# a_n803_n800# a_1519_n800# a_n2093_n800#
+ a_803_n855# a_n2035_n855#
X0 a_n1577_n800# a_n1777_n855# a_n1835_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X1 a_1519_n800# a_1319_n855# a_1261_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X2 a_n1061_n800# a_n1261_n855# a_n1319_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X3 a_745_n800# a_545_n855# a_487_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X4 a_1003_n800# a_803_n855# a_745_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X5 a_487_n800# a_287_n855# a_229_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X6 a_2035_n800# a_1835_n855# a_1777_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X7 a_1777_n800# a_1577_n855# a_1519_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X8 a_1261_n800# a_1061_n855# a_1003_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X9 a_n1835_n800# a_n2035_n855# a_n2093_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X10 a_n2093_n800# a_n2293_n855# a_n2351_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=1
X11 a_n29_n800# a_n229_n855# a_n287_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X12 a_229_n800# a_29_n855# a_n29_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X13 a_n1319_n800# a_n1519_n855# a_n1577_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X14 a_n545_n800# a_n745_n855# a_n803_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X15 a_2293_n800# a_2093_n855# a_2035_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=1
X16 a_n803_n800# a_n1003_n855# a_n1061_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X17 a_n287_n800# a_n487_n855# a_n545_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_79TVLH a_3067_n300# a_1777_n300# a_n2609_n300#
+ a_1061_n355# a_n2293_n355# a_n2351_n300# a_229_n300# a_n1577_n300# a_n1519_n355#
+ a_2035_n300# a_n487_n355# a_n545_n300# a_n1261_n355# a_2609_n355# a_545_n355# a_n3517_n522#
+ a_2351_n355# a_1003_n300# a_1577_n355# a_n2867_n300# a_n2809_n355# a_3325_n300#
+ a_n2551_n355# a_487_n300# a_n29_n300# a_n3067_n355# a_29_n355# a_n1777_n355# a_2293_n300#
+ a_n1835_n300# a_n3125_n300# a_n745_n355# a_2867_n355# a_1519_n300# a_n803_n300#
+ a_n2093_n300# a_803_n355# a_n2035_n355# a_1261_n300# a_n1319_n300# a_3125_n355#
+ a_1835_n355# a_n287_n300# a_n229_n355# a_n1061_n300# a_287_n355# a_n1003_n355# a_2809_n300#
+ a_745_n300# a_2093_n355# a_n3383_n300# a_n3325_n355# a_2551_n300# a_1319_n355#
X0 a_2809_n300# a_2609_n355# a_2551_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1 a_n2351_n300# a_n2551_n355# a_n2609_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X2 a_n2093_n300# a_n2293_n355# a_n2351_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X3 a_229_n300# a_29_n355# a_n29_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X4 a_n29_n300# a_n229_n355# a_n287_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X5 a_3067_n300# a_2867_n355# a_2809_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X6 a_n1319_n300# a_n1519_n355# a_n1577_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X7 a_n545_n300# a_n745_n355# a_n803_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X8 a_2293_n300# a_2093_n355# a_2035_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X9 a_2551_n300# a_2351_n355# a_2293_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X10 a_n3125_n300# a_n3325_n355# a_n3383_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X11 a_n2867_n300# a_n3067_n355# a_n3125_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X12 a_n803_n300# a_n1003_n355# a_n1061_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X13 a_n287_n300# a_n487_n355# a_n545_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X14 a_n1577_n300# a_n1777_n355# a_n1835_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X15 a_1519_n300# a_1319_n355# a_1261_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X16 a_3325_n300# a_3125_n355# a_3067_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X17 a_n1061_n300# a_n1261_n355# a_n1319_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X18 a_1003_n300# a_803_n355# a_745_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X19 a_487_n300# a_287_n355# a_229_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X20 a_745_n300# a_545_n355# a_487_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X21 a_2035_n300# a_1835_n355# a_1777_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X22 a_n2609_n300# a_n2809_n355# a_n2867_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X23 a_1777_n300# a_1577_n355# a_1519_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X24 a_1261_n300# a_1061_n355# a_1003_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X25 a_n1835_n300# a_n2035_n355# a_n2093_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_U73S5M a_229_n1000# a_n803_n1000# a_545_n1055#
+ a_29_n1055# a_n487_n1055# a_n4549_n1222# a_n3641_n1000# a_3841_n1000# a_3067_n1000#
+ a_3383_n1055# a_2867_n1055# a_2551_n1000# a_n2351_n1000# a_n1835_n1000# a_n4415_n1000#
+ a_2093_n1055# a_n4099_n1055# a_1577_n1055# a_803_n1055# a_n745_n1055# a_n1003_n1055#
+ a_n1061_n1000# a_4157_n1055# a_n3583_n1055# a_1261_n1000# a_n3125_n1000# a_3641_n1055#
+ a_3325_n1000# a_2809_n1000# a_n2609_n1000# a_n2293_n1055# a_n1777_n1055# a_2035_n1000#
+ a_2351_n1055# a_n4357_n1055# a_1519_n1000# a_n1319_n1000# a_n3899_n1000# a_1835_n1055#
+ a_487_n1000# a_n229_n1055# a_n3841_n1055# a_n287_n1000# a_1061_n1055# a_n3067_n1055#
+ a_3125_n1055# a_n2551_n1055# a_2609_n1055# a_1319_n1055# a_n1261_n1055# a_4099_n1000#
+ a_745_n1000# a_3899_n1055# a_1003_n1000# a_n545_n1000# a_287_n1055# a_n2809_n1055#
+ a_n3325_n1055# a_3583_n1000# a_n3383_n1000# a_n2867_n1000# a_n2035_n1055# a_n2093_n1000#
+ a_n1519_n1055# a_2293_n1000# a_n1577_n1000# a_4357_n1000# a_1777_n1000# a_n29_n1000#
+ a_n4157_n1000#
X0 a_3067_n1000# a_2867_n1055# a_2809_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X1 a_n1319_n1000# a_n1519_n1055# a_n1577_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X2 a_n545_n1000# a_n745_n1055# a_n803_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X3 a_2293_n1000# a_2093_n1055# a_2035_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X4 a_2551_n1000# a_2351_n1055# a_2293_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X5 a_n3125_n1000# a_n3325_n1055# a_n3383_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X6 a_n2867_n1000# a_n3067_n1055# a_n3125_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X7 a_n803_n1000# a_n1003_n1055# a_n1061_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X8 a_n287_n1000# a_n487_n1055# a_n545_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X9 a_n3641_n1000# a_n3841_n1055# a_n3899_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X10 a_n1577_n1000# a_n1777_n1055# a_n1835_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X11 a_1519_n1000# a_1319_n1055# a_1261_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X12 a_n3383_n1000# a_n3583_n1055# a_n3641_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X13 a_3325_n1000# a_3125_n1055# a_3067_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X14 a_n1061_n1000# a_n1261_n1055# a_n1319_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X15 a_745_n1000# a_545_n1055# a_487_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X16 a_1003_n1000# a_803_n1055# a_745_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X17 a_487_n1000# a_287_n1055# a_229_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X18 a_2035_n1000# a_1835_n1055# a_1777_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X19 a_4099_n1000# a_3899_n1055# a_3841_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X20 a_n2609_n1000# a_n2809_n1055# a_n2867_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X21 a_1777_n1000# a_1577_n1055# a_1519_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X22 a_3841_n1000# a_3641_n1055# a_3583_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X23 a_1261_n1000# a_1061_n1055# a_1003_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X24 a_3583_n1000# a_3383_n1055# a_3325_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X25 a_n4157_n1000# a_n4357_n1055# a_n4415_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=1
X26 a_n3899_n1000# a_n4099_n1055# a_n4157_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X27 a_n1835_n1000# a_n2035_n1055# a_n2093_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X28 a_2809_n1000# a_2609_n1055# a_2551_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X29 a_n2351_n1000# a_n2551_n1055# a_n2609_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X30 a_4357_n1000# a_4157_n1055# a_4099_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=1
X31 a_n2093_n1000# a_n2293_n1055# a_n2351_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X32 a_n29_n1000# a_n229_n1055# a_n287_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X33 a_229_n1000# a_29_n1055# a_n29_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_PP2RNK a_29_n964# a_n2351_n900# a_229_n900# a_2867_n964#
+ a_n745_n964# a_n1577_n900# a_2035_n900# a_803_n964# a_n2035_n964# a_n545_n900# w_n3325_n1197#
+ a_1835_n964# a_1003_n900# a_n229_n964# a_n1003_n964# a_287_n964# a_n2867_n900# a_2093_n964#
+ a_487_n900# a_n29_n900# a_2293_n900# a_n3125_n900# a_1319_n964# a_n1835_n900# a_1061_n964#
+ a_n2293_n964# a_n803_n900# a_1519_n900# a_n2093_n900# a_n1519_n964# a_1261_n900#
+ a_n487_n964# a_n1261_n964# a_2609_n964# a_n1319_n900# a_545_n964# a_n287_n900# a_2351_n964#
+ a_n1061_n900# a_1577_n964# a_2809_n900# a_745_n900# a_n2809_n964# a_2551_n900# a_n2551_n964#
+ a_3067_n900# a_1777_n900# a_n2609_n900# a_n1777_n964# a_n3067_n964#
X0 a_1261_n900# a_1061_n964# a_1003_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1 a_n1835_n900# a_n2035_n964# a_n2093_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X2 a_2809_n900# a_2609_n964# a_2551_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X3 a_n2351_n900# a_n2551_n964# a_n2609_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X4 a_n2093_n900# a_n2293_n964# a_n2351_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X5 a_n29_n900# a_n229_n964# a_n287_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X6 a_229_n900# a_29_n964# a_n29_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X7 a_3067_n900# a_2867_n964# a_2809_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X8 a_2551_n900# a_2351_n964# a_2293_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X9 a_n1319_n900# a_n1519_n964# a_n1577_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X10 a_n545_n900# a_n745_n964# a_n803_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X11 a_2293_n900# a_2093_n964# a_2035_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X12 a_n2867_n900# a_n3067_n964# a_n3125_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X13 a_n803_n900# a_n1003_n964# a_n1061_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X14 a_n287_n900# a_n487_n964# a_n545_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X15 a_n1577_n900# a_n1777_n964# a_n1835_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X16 a_1519_n900# a_1319_n964# a_1261_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X17 a_n1061_n900# a_n1261_n964# a_n1319_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X18 a_745_n900# a_545_n964# a_487_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X19 a_1003_n900# a_803_n964# a_745_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X20 a_487_n900# a_287_n964# a_229_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X21 a_2035_n900# a_1835_n964# a_1777_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X22 a_n2609_n900# a_n2809_n964# a_n2867_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X23 a_1777_n900# a_1577_n964# a_1519_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QTY6H6 a_1261_n200# a_n487_n264# a_n1261_n264#
+ a_n1319_n200# a_545_n264# a_n287_n200# a_n1061_n200# a_745_n200# a_29_n264# a_229_n200#
+ a_n745_n264# a_n1577_n200# a_803_n264# a_n545_n200# a_1003_n200# a_n229_n264# a_n1003_n264#
+ a_287_n264# a_487_n200# a_n29_n200# a_1319_n264# a_1061_n264# w_n1777_n497# a_n803_n200#
+ a_1519_n200# a_n1519_n264#
X0 a_487_n200# a_287_n264# a_229_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_1261_n200# a_1061_n264# a_1003_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_n29_n200# a_n229_n264# a_n287_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_229_n200# a_29_n264# a_n29_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_n1319_n200# a_n1519_n264# a_n1577_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X5 a_n545_n200# a_n745_n264# a_n803_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_n803_n200# a_n1003_n264# a_n1061_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_n287_n200# a_n487_n264# a_n545_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_1519_n200# a_1319_n264# a_1261_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X9 a_n1061_n200# a_n1261_n264# a_n1319_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_745_n200# a_545_n264# a_487_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_1003_n200# a_803_n264# a_745_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NT3TPY a_n287_n255# a_n345_n200# a_345_n255#
+ a_n445_n255# a_129_n200# a_n503_n200# a_287_n200# a_445_n200# a_n637_n422# a_n29_n200#
+ a_29_n255# a_n187_n200# a_n129_n255# a_187_n255#
X0 a_n187_n200# a_n287_n255# a_n345_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X1 a_287_n200# a_187_n255# a_129_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X2 a_n345_n200# a_n445_n255# a_n503_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X3 a_129_n200# a_29_n255# a_n29_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X4 a_445_n200# a_345_n255# a_287_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X5 a_n29_n200# a_n129_n255# a_n187_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_5X2ZTR a_n2093_n200# a_803_n255# a_n2035_n255#
+ a_n3841_n255# a_n5131_n255# a_1261_n200# a_n4357_n255# a_3583_n200# a_n1319_n200#
+ a_n4415_n200# a_4931_n255# a_3125_n255# a_1835_n255# a_n287_n200# a_n229_n255# a_4099_n200#
+ a_n1061_n200# a_287_n255# a_n1003_n255# a_2809_n200# a_745_n200# a_n3383_n200# a_2093_n255#
+ a_n3325_n255# a_2551_n200# a_3067_n200# a_4415_n255# a_1319_n255# a_4873_n200# a_1777_n200#
+ a_n2609_n200# a_n2293_n255# a_1061_n255# a_n5323_n422# a_n2351_n200# a_229_n200#
+ a_3383_n255# a_n1577_n200# a_n4673_n200# a_n1519_n255# a_n4615_n255# a_5131_n200#
+ a_3841_n200# a_2035_n200# a_n487_n255# a_n545_n200# a_n3899_n200# a_n5189_n200#
+ a_n1261_n255# a_4357_n200# a_2609_n255# a_545_n255# a_n3583_n255# a_n3641_n200#
+ a_2351_n255# a_1003_n200# a_n4099_n255# a_n4157_n200# a_4673_n255# a_1577_n255#
+ a_3325_n200# a_n2867_n200# a_n2809_n255# a_3899_n255# a_n2551_n255# a_487_n200#
+ a_n29_n200# a_n3067_n255# a_2293_n200# a_29_n255# a_n1777_n255# a_n4873_n255# a_n1835_n200#
+ a_n3125_n200# a_n4931_n200# a_3641_n255# a_4157_n255# a_n745_n255# a_n803_n200#
+ a_2867_n255# a_4615_n200# a_1519_n200#
X0 a_2035_n200# a_1835_n255# a_1777_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_4099_n200# a_3899_n255# a_3841_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_n2609_n200# a_n2809_n255# a_n2867_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_1777_n200# a_1577_n255# a_1519_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_3841_n200# a_3641_n255# a_3583_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_n4415_n200# a_n4615_n255# a_n4673_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_1261_n200# a_1061_n255# a_1003_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_3583_n200# a_3383_n255# a_3325_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_n4157_n200# a_n4357_n255# a_n4415_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_n3899_n200# a_n4099_n255# a_n4157_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_n1835_n200# a_n2035_n255# a_n2093_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_n4673_n200# a_n4873_n255# a_n4931_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X12 a_2809_n200# a_2609_n255# a_2551_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X13 a_n2351_n200# a_n2551_n255# a_n2609_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X14 a_4357_n200# a_4157_n255# a_4099_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X15 a_4615_n200# a_4415_n255# a_4357_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X16 a_n2093_n200# a_n2293_n255# a_n2351_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X17 a_n29_n200# a_n229_n255# a_n287_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X18 a_229_n200# a_29_n255# a_n29_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X19 a_3067_n200# a_2867_n255# a_2809_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X20 a_5131_n200# a_4931_n255# a_4873_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X21 a_4873_n200# a_4673_n255# a_4615_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X22 a_n1319_n200# a_n1519_n255# a_n1577_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X23 a_n545_n200# a_n745_n255# a_n803_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X24 a_2293_n200# a_2093_n255# a_2035_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X25 a_2551_n200# a_2351_n255# a_2293_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X26 a_n3125_n200# a_n3325_n255# a_n3383_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X27 a_n2867_n200# a_n3067_n255# a_n3125_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X28 a_n803_n200# a_n1003_n255# a_n1061_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X29 a_n287_n200# a_n487_n255# a_n545_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X30 a_n4931_n200# a_n5131_n255# a_n5189_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X31 a_n3641_n200# a_n3841_n255# a_n3899_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X32 a_n1577_n200# a_n1777_n255# a_n1835_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X33 a_1519_n200# a_1319_n255# a_1261_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X34 a_n3383_n200# a_n3583_n255# a_n3641_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X35 a_3325_n200# a_3125_n255# a_3067_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X36 a_n1061_n200# a_n1261_n255# a_n1319_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X37 a_745_n200# a_545_n255# a_487_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X38 a_1003_n200# a_803_n255# a_745_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X39 a_487_n200# a_287_n255# a_229_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WK95DB a_n819_n450# a_n345_n450# a_29_n505# a_n129_n505#
+ a_187_n505# a_129_n450# a_n503_n450# a_n287_n505# a_345_n505# a_287_n450# a_n661_n450#
+ a_n445_n505# a_503_n505# a_445_n450# a_n603_n505# a_661_n505# a_603_n450# a_n761_n505#
+ a_761_n450# a_n953_n672# a_n29_n450# a_n187_n450#
X0 a_129_n450# a_29_n505# a_n29_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X1 a_445_n450# a_345_n505# a_287_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X2 a_n503_n450# a_n603_n505# a_n661_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X3 a_n29_n450# a_n129_n505# a_n187_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X4 a_603_n450# a_503_n505# a_445_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X5 a_n661_n450# a_n761_n505# a_n819_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=0.5
X6 a_n187_n450# a_n287_n505# a_n345_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X7 a_761_n450# a_661_n505# a_603_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=0.5
X8 a_287_n450# a_187_n505# a_129_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X9 a_n345_n450# a_n445_n505# a_n503_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PGZBW9 a_1061_n655# a_n2293_n655# a_n2351_n600#
+ a_229_n600# a_n1577_n600# a_n1519_n655# a_2035_n600# a_n487_n655# a_n1261_n655#
+ a_n545_n600# a_2609_n655# a_545_n655# a_2351_n655# a_n3517_n822# a_1003_n600# a_1577_n655#
+ a_n2867_n600# a_n2809_n655# a_3325_n600# a_n2551_n655# a_n29_n600# a_487_n600# a_n1777_n655#
+ a_n3067_n655# a_2293_n600# a_n3125_n600# a_29_n655# a_n1835_n600# a_2867_n655# a_n745_n655#
+ a_n803_n600# a_1519_n600# a_n2093_n600# a_803_n655# a_n2035_n655# a_1261_n600# a_3125_n655#
+ a_n1319_n600# a_1835_n655# a_n287_n600# a_n1061_n600# a_n229_n655# a_n1003_n655#
+ a_287_n655# a_2809_n600# a_2093_n655# a_745_n600# a_n3383_n600# a_n3325_n655# a_2551_n600#
+ a_3067_n600# a_1777_n600# a_n2609_n600# a_1319_n655#
X0 a_2809_n600# a_2609_n655# a_2551_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X1 a_n2351_n600# a_n2551_n655# a_n2609_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X2 a_n2093_n600# a_n2293_n655# a_n2351_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X3 a_n29_n600# a_n229_n655# a_n287_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X4 a_229_n600# a_29_n655# a_n29_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X5 a_3067_n600# a_2867_n655# a_2809_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X6 a_n1319_n600# a_n1519_n655# a_n1577_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X7 a_2551_n600# a_2351_n655# a_2293_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X8 a_n3125_n600# a_n3325_n655# a_n3383_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=1
X9 a_n545_n600# a_n745_n655# a_n803_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X10 a_n287_n600# a_n487_n655# a_n545_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X11 a_2293_n600# a_2093_n655# a_2035_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X12 a_n2867_n600# a_n3067_n655# a_n3125_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X13 a_n803_n600# a_n1003_n655# a_n1061_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X14 a_n1577_n600# a_n1777_n655# a_n1835_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X15 a_1519_n600# a_1319_n655# a_1261_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X16 a_n1061_n600# a_n1261_n655# a_n1319_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X17 a_3325_n600# a_3125_n655# a_3067_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=1
X18 a_1003_n600# a_803_n655# a_745_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X19 a_745_n600# a_545_n655# a_487_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X20 a_487_n600# a_287_n655# a_229_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X21 a_1777_n600# a_1577_n655# a_1519_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X22 a_2035_n600# a_1835_n655# a_1777_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X23 a_n2609_n600# a_n2809_n655# a_n2867_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X24 a_1261_n600# a_1061_n655# a_1003_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X25 a_n1835_n600# a_n2035_n655# a_n2093_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3QL9S5 a_n50_n497# a_50_n400# w_n308_n697# a_n108_n400#
X0 a_50_n400# a_n50_n497# a_n108_n400# w_n308_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_U4Z9ZD a_761_n400# a_503_n464# a_n29_n400# a_n603_n464#
+ a_661_n464# a_n187_n400# a_n761_n464# a_n819_n400# a_n345_n400# a_129_n400# a_n503_n400#
+ w_n1019_n697# a_287_n400# a_n661_n400# a_29_n464# a_n129_n464# a_187_n464# a_445_n400#
+ a_n287_n464# a_345_n464# a_603_n400# a_n445_n464#
X0 a_n503_n400# a_n603_n464# a_n661_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X1 a_n29_n400# a_n129_n464# a_n187_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 a_603_n400# a_503_n464# a_445_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n661_n400# a_n761_n464# a_n819_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X4 a_n187_n400# a_n287_n464# a_n345_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X5 a_761_n400# a_661_n464# a_603_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X6 a_287_n400# a_187_n464# a_129_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X7 a_n345_n400# a_n445_n464# a_n503_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X8 a_129_n400# a_29_n464# a_n29_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X9 a_445_n400# a_345_n464# a_287_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QSKB8C a_287_n464# a_n1003_n464# a_n2867_n400#
+ a_n4157_n400# a_2093_n464# a_3325_n400# a_n3325_n464# a_487_n400# a_n29_n400# a_4415_n464#
+ a_1319_n464# a_2293_n400# a_n1835_n400# a_n3125_n400# a_n2293_n464# a_n4931_n400#
+ a_1061_n464# a_1519_n400# a_n803_n400# a_3383_n464# a_4615_n400# a_n2093_n400# a_n1519_n464#
+ a_n4615_n464# a_1261_n400# a_n487_n464# a_n1261_n464# w_n5131_n697# a_n1319_n400#
+ a_2609_n464# a_545_n464# a_3583_n400# a_n287_n400# a_n4415_n400# a_n3583_n464# a_4099_n400#
+ a_n1061_n400# a_2351_n464# a_n4099_n464# a_2809_n400# a_4673_n464# a_1577_n464#
+ a_745_n400# a_n3383_n400# a_n2809_n464# a_2551_n400# a_3899_n464# a_n2551_n464#
+ a_4873_n400# a_3067_n400# a_1777_n400# a_n2609_n400# a_n3067_n464# a_3641_n464#
+ a_29_n464# a_n1777_n464# a_n4873_n464# a_n2351_n400# a_4157_n464# a_n745_n464# a_229_n400#
+ a_n1577_n400# a_n4673_n400# a_2867_n464# a_2035_n400# a_803_n464# a_n2035_n464#
+ a_3841_n400# a_n3841_n464# a_4357_n400# a_n545_n400# a_n3899_n400# a_3125_n464#
+ a_n4357_n464# a_1835_n464# a_1003_n400# a_n3641_n400# a_n229_n464#
X0 a_4873_n400# a_4673_n464# a_4615_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X1 a_n1319_n400# a_n1519_n464# a_n1577_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X2 a_n545_n400# a_n745_n464# a_n803_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 a_2293_n400# a_2093_n464# a_2035_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X4 a_2551_n400# a_2351_n464# a_2293_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X5 a_n3125_n400# a_n3325_n464# a_n3383_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X6 a_n2867_n400# a_n3067_n464# a_n3125_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X7 a_n803_n400# a_n1003_n464# a_n1061_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X8 a_n287_n400# a_n487_n464# a_n545_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X9 a_n3641_n400# a_n3841_n464# a_n3899_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X10 a_n1577_n400# a_n1777_n464# a_n1835_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X11 a_n3383_n400# a_n3583_n464# a_n3641_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X12 a_1519_n400# a_1319_n464# a_1261_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X13 a_3325_n400# a_3125_n464# a_3067_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X14 a_n1061_n400# a_n1261_n464# a_n1319_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X15 a_1003_n400# a_803_n464# a_745_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X16 a_487_n400# a_287_n464# a_229_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X17 a_745_n400# a_545_n464# a_487_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X18 a_2035_n400# a_1835_n464# a_1777_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X19 a_4099_n400# a_3899_n464# a_3841_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X20 a_n2609_n400# a_n2809_n464# a_n2867_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X21 a_1777_n400# a_1577_n464# a_1519_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X22 a_3841_n400# a_3641_n464# a_3583_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X23 a_n4415_n400# a_n4615_n464# a_n4673_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X24 a_1261_n400# a_1061_n464# a_1003_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X25 a_3583_n400# a_3383_n464# a_3325_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X26 a_n4157_n400# a_n4357_n464# a_n4415_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X27 a_n3899_n400# a_n4099_n464# a_n4157_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X28 a_n1835_n400# a_n2035_n464# a_n2093_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X29 a_n4673_n400# a_n4873_n464# a_n4931_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X30 a_2809_n400# a_2609_n464# a_2551_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X31 a_n2351_n400# a_n2551_n464# a_n2609_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X32 a_4357_n400# a_4157_n464# a_4099_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X33 a_4615_n400# a_4415_n464# a_4357_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X34 a_n2093_n400# a_n2293_n464# a_n2351_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X35 a_229_n400# a_29_n464# a_n29_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X36 a_n29_n400# a_n229_n464# a_n287_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X37 a_3067_n400# a_2867_n464# a_2809_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QRKB8C a_287_n464# a_n1003_n464# a_n2867_n400#
+ a_n4157_n400# a_2093_n464# a_3325_n400# a_n3325_n464# a_487_n400# a_n29_n400# a_4415_n464#
+ a_1319_n464# a_2293_n400# a_n1835_n400# a_n3125_n400# a_n2293_n464# a_1061_n464#
+ w_n4873_n697# a_1519_n400# a_n803_n400# a_3383_n464# a_4615_n400# a_n2093_n400#
+ a_n1519_n464# a_n4615_n464# a_1261_n400# a_n487_n464# a_n1261_n464# a_n1319_n400#
+ a_2609_n464# a_545_n464# a_3583_n400# a_n287_n400# a_n4415_n400# a_n3583_n464# a_4099_n400#
+ a_n1061_n400# a_2351_n464# a_n4099_n464# a_2809_n400# a_1577_n464# a_745_n400# a_n3383_n400#
+ a_n2809_n464# a_2551_n400# a_3899_n464# a_n2551_n464# a_3067_n400# a_1777_n400#
+ a_n2609_n400# a_n3067_n464# a_3641_n464# a_29_n464# a_n1777_n464# a_n2351_n400#
+ a_4157_n464# a_n745_n464# a_229_n400# a_n1577_n400# a_n4673_n400# a_2867_n464# a_2035_n400#
+ a_803_n464# a_n2035_n464# a_3841_n400# a_n3841_n464# a_4357_n400# a_n545_n400# a_n3899_n400#
+ a_3125_n464# a_n4357_n464# a_1835_n464# a_1003_n400# a_n3641_n400# a_n229_n464#
X0 a_n1319_n400# a_n1519_n464# a_n1577_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X1 a_n545_n400# a_n745_n464# a_n803_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X2 a_2293_n400# a_2093_n464# a_2035_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 a_2551_n400# a_2351_n464# a_2293_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X4 a_n3125_n400# a_n3325_n464# a_n3383_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X5 a_n2867_n400# a_n3067_n464# a_n3125_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X6 a_n803_n400# a_n1003_n464# a_n1061_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X7 a_n287_n400# a_n487_n464# a_n545_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X8 a_n3641_n400# a_n3841_n464# a_n3899_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X9 a_n1577_n400# a_n1777_n464# a_n1835_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X10 a_n3383_n400# a_n3583_n464# a_n3641_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X11 a_1519_n400# a_1319_n464# a_1261_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X12 a_3325_n400# a_3125_n464# a_3067_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X13 a_n1061_n400# a_n1261_n464# a_n1319_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X14 a_1003_n400# a_803_n464# a_745_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X15 a_487_n400# a_287_n464# a_229_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X16 a_745_n400# a_545_n464# a_487_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X17 a_2035_n400# a_1835_n464# a_1777_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X18 a_4099_n400# a_3899_n464# a_3841_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X19 a_n2609_n400# a_n2809_n464# a_n2867_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X20 a_1777_n400# a_1577_n464# a_1519_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X21 a_3841_n400# a_3641_n464# a_3583_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X22 a_n4415_n400# a_n4615_n464# a_n4673_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X23 a_1261_n400# a_1061_n464# a_1003_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X24 a_3583_n400# a_3383_n464# a_3325_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X25 a_n4157_n400# a_n4357_n464# a_n4415_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X26 a_n3899_n400# a_n4099_n464# a_n4157_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X27 a_n1835_n400# a_n2035_n464# a_n2093_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X28 a_2809_n400# a_2609_n464# a_2551_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X29 a_n2351_n400# a_n2551_n464# a_n2609_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X30 a_4357_n400# a_4157_n464# a_4099_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X31 a_4615_n400# a_4415_n464# a_4357_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X32 a_n2093_n400# a_n2293_n464# a_n2351_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X33 a_229_n400# a_29_n464# a_n29_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X34 a_n29_n400# a_n229_n464# a_n287_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X35 a_3067_n400# a_2867_n464# a_2809_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_EVM3FM a_29_n964# a_n129_n964# a_187_n964# a_445_n900#
+ a_n287_n964# a_345_n964# a_603_n900# a_n445_n964# a_761_n900# a_503_n964# a_n29_n900#
+ a_n603_n964# a_661_n964# a_n187_n900# a_n761_n964# a_n819_n900# a_n345_n900# a_129_n900#
+ a_n503_n900# w_n1019_n1197# a_n661_n900# a_287_n900#
X0 a_n187_n900# a_n287_n964# a_n345_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X1 a_761_n900# a_661_n964# a_603_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=0.5
X2 a_287_n900# a_187_n964# a_129_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X3 a_n345_n900# a_n445_n964# a_n503_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X4 a_129_n900# a_29_n964# a_n29_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X5 a_445_n900# a_345_n964# a_287_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X6 a_n503_n900# a_n603_n964# a_n661_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X7 a_n29_n900# a_n129_n964# a_n187_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X8 a_603_n900# a_503_n964# a_445_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X9 a_n661_n900# a_n761_n964# a_n819_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DL2ZHN a_n2093_n200# a_803_n255# a_n2035_n255#
+ a_n3841_n255# a_1261_n200# a_n4357_n255# a_3583_n200# a_n1319_n200# a_n4415_n200#
+ a_3125_n255# a_1835_n255# a_n287_n200# a_n229_n255# a_4099_n200# a_n1061_n200# a_287_n255#
+ a_n1003_n255# a_2809_n200# a_745_n200# a_n3383_n200# a_2093_n255# a_n3325_n255#
+ a_2551_n200# a_3067_n200# a_4415_n255# a_1319_n255# a_4873_n200# a_1777_n200# a_n2609_n200#
+ a_n2293_n255# a_1061_n255# a_n2351_n200# a_229_n200# a_3383_n255# a_n1577_n200#
+ a_n4673_n200# a_n1519_n255# a_n4615_n255# a_3841_n200# a_2035_n200# a_n487_n255#
+ a_n545_n200# a_n3899_n200# a_n1261_n255# a_4357_n200# a_2609_n255# a_545_n255# a_n3583_n255#
+ a_n3641_n200# a_2351_n255# a_1003_n200# a_n4099_n255# a_n4157_n200# a_4673_n255#
+ a_1577_n255# a_3325_n200# a_n2867_n200# a_n2809_n255# a_3899_n255# a_n2551_n255#
+ a_487_n200# a_n29_n200# a_n3067_n255# a_2293_n200# a_29_n255# a_n1777_n255# a_n4873_n255#
+ a_n1835_n200# a_n3125_n200# a_n4931_n200# a_3641_n255# a_4157_n255# a_n745_n255#
+ a_n803_n200# a_2867_n255# a_4615_n200# a_1519_n200# a_n5065_n422#
X0 a_2035_n200# a_1835_n255# a_1777_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_4099_n200# a_3899_n255# a_3841_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_n2609_n200# a_n2809_n255# a_n2867_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_1777_n200# a_1577_n255# a_1519_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_3841_n200# a_3641_n255# a_3583_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_n4415_n200# a_n4615_n255# a_n4673_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_1261_n200# a_1061_n255# a_1003_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_3583_n200# a_3383_n255# a_3325_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_n4157_n200# a_n4357_n255# a_n4415_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_n3899_n200# a_n4099_n255# a_n4157_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_n1835_n200# a_n2035_n255# a_n2093_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_n4673_n200# a_n4873_n255# a_n4931_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X12 a_2809_n200# a_2609_n255# a_2551_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X13 a_n2351_n200# a_n2551_n255# a_n2609_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X14 a_4357_n200# a_4157_n255# a_4099_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X15 a_4615_n200# a_4415_n255# a_4357_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X16 a_n2093_n200# a_n2293_n255# a_n2351_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X17 a_n29_n200# a_n229_n255# a_n287_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X18 a_229_n200# a_29_n255# a_n29_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X19 a_3067_n200# a_2867_n255# a_2809_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X20 a_4873_n200# a_4673_n255# a_4615_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X21 a_n1319_n200# a_n1519_n255# a_n1577_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X22 a_n545_n200# a_n745_n255# a_n803_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X23 a_2293_n200# a_2093_n255# a_2035_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X24 a_2551_n200# a_2351_n255# a_2293_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X25 a_n3125_n200# a_n3325_n255# a_n3383_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X26 a_n2867_n200# a_n3067_n255# a_n3125_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X27 a_n803_n200# a_n1003_n255# a_n1061_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X28 a_n287_n200# a_n487_n255# a_n545_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X29 a_n3641_n200# a_n3841_n255# a_n3899_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X30 a_n1577_n200# a_n1777_n255# a_n1835_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X31 a_1519_n200# a_1319_n255# a_1261_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X32 a_n3383_n200# a_n3583_n255# a_n3641_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X33 a_3325_n200# a_3125_n255# a_3067_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X34 a_n1061_n200# a_n1261_n255# a_n1319_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X35 a_745_n200# a_545_n255# a_487_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X36 a_1003_n200# a_803_n255# a_745_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X37 a_487_n200# a_287_n255# a_229_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_HG2LSW a_n100_n205# a_100_n150# a_n292_n372#
+ a_n158_n150#
X0 a_100_n150# a_n100_n205# a_n158_n150# a_n292_n372# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_N64HU4 a_3235_n255# a_n1861_n200# a_n1803_n255#
+ a_n3827_n422# a_n2777_n200# a_n1345_n255# a_n2719_n255# a_3635_n200# a_2261_n200#
+ a_n1403_n200# a_3177_n200# a_n2319_n200# a_1861_n255# a_2777_n255# a_1403_n255#
+ a_n887_n255# a_n945_n200# a_945_n255# a_2319_n255# a_n487_n200# a_n429_n255# a_1803_n200#
+ a_487_n255# a_2719_n200# a_1345_n200# a_n29_n200# a_n3693_n200# a_n2261_n255# a_n3635_n255#
+ a_887_n200# a_29_n255# a_n3177_n255# a_n3235_n200# a_429_n200#
X0 a_n2319_n200# a_n2719_n255# a_n2777_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X1 a_n2777_n200# a_n3177_n255# a_n3235_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X2 a_2261_n200# a_1861_n255# a_1803_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X3 a_n945_n200# a_n1345_n255# a_n1403_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X4 a_3635_n200# a_3235_n255# a_3177_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=2
X5 a_429_n200# a_29_n255# a_n29_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X6 a_1803_n200# a_1403_n255# a_1345_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X7 a_887_n200# a_487_n255# a_429_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X8 a_3177_n200# a_2777_n255# a_2719_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X9 a_n3235_n200# a_n3635_n255# a_n3693_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=2
X10 a_n487_n200# a_n887_n255# a_n945_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X11 a_n1403_n200# a_n1803_n255# a_n1861_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X12 a_2719_n200# a_2319_n255# a_2261_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X13 a_n1861_n200# a_n2261_n255# a_n2319_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X14 a_n29_n200# a_n429_n255# a_n487_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X15 a_1345_n200# a_945_n255# a_887_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UGZTXE a_1061_n655# a_n2293_n655# a_n2351_n600#
+ a_229_n600# a_n1577_n600# a_3383_n655# a_n1519_n655# a_2035_n600# a_n487_n655# a_n1261_n655#
+ a_n545_n600# a_2609_n655# a_545_n655# a_2351_n655# a_n3583_n655# a_1003_n600# a_n3641_n600#
+ a_1577_n655# a_n2867_n600# a_n2809_n655# a_3325_n600# a_n2551_n655# a_n29_n600#
+ a_487_n600# a_n1777_n655# a_n3067_n655# a_2293_n600# a_n3125_n600# a_29_n655# a_n1835_n600#
+ a_2867_n655# a_n745_n655# a_n803_n600# a_1519_n600# a_n2093_n600# a_803_n655# a_n2035_n655#
+ a_n3775_n822# a_1261_n600# a_3125_n655# a_3583_n600# a_n1319_n600# a_1835_n655#
+ a_n287_n600# a_n1061_n600# a_n229_n655# a_n1003_n655# a_287_n655# a_2809_n600# a_2093_n655#
+ a_745_n600# a_n3383_n600# a_n3325_n655# a_2551_n600# a_3067_n600# a_1777_n600# a_n2609_n600#
+ a_1319_n655#
X0 a_2809_n600# a_2609_n655# a_2551_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X1 a_n2351_n600# a_n2551_n655# a_n2609_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X2 a_n2093_n600# a_n2293_n655# a_n2351_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X3 a_n29_n600# a_n229_n655# a_n287_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X4 a_229_n600# a_29_n655# a_n29_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X5 a_3067_n600# a_2867_n655# a_2809_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X6 a_n1319_n600# a_n1519_n655# a_n1577_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X7 a_2551_n600# a_2351_n655# a_2293_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X8 a_n3125_n600# a_n3325_n655# a_n3383_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X9 a_n545_n600# a_n745_n655# a_n803_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X10 a_n287_n600# a_n487_n655# a_n545_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X11 a_2293_n600# a_2093_n655# a_2035_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X12 a_n2867_n600# a_n3067_n655# a_n3125_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X13 a_n803_n600# a_n1003_n655# a_n1061_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X14 a_n1577_n600# a_n1777_n655# a_n1835_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X15 a_1519_n600# a_1319_n655# a_1261_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X16 a_n3383_n600# a_n3583_n655# a_n3641_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=1
X17 a_n1061_n600# a_n1261_n655# a_n1319_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X18 a_3325_n600# a_3125_n655# a_3067_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X19 a_1003_n600# a_803_n655# a_745_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X20 a_745_n600# a_545_n655# a_487_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X21 a_487_n600# a_287_n655# a_229_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X22 a_1777_n600# a_1577_n655# a_1519_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X23 a_2035_n600# a_1835_n655# a_1777_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X24 a_n2609_n600# a_n2809_n655# a_n2867_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X25 a_3583_n600# a_3383_n655# a_3325_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=1
X26 a_1261_n600# a_1061_n655# a_1003_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X27 a_n1835_n600# a_n2035_n655# a_n2093_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Q46EE6 a_1261_n200# a_n487_n264# a_n1261_n264#
+ w_n2035_n497# a_n1319_n200# a_545_n264# a_n287_n200# a_n1061_n200# a_1577_n264#
+ a_745_n200# a_1777_n200# a_n1777_n264# a_29_n264# a_229_n200# a_n745_n264# a_n1577_n200#
+ a_803_n264# a_n545_n200# a_1003_n200# a_n229_n264# a_n1003_n264# a_287_n264# a_487_n200#
+ a_n29_n200# a_1319_n264# a_n1835_n200# a_1061_n264# a_n803_n200# a_1519_n200# a_n1519_n264#
X0 a_487_n200# a_287_n264# a_229_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_1777_n200# a_1577_n264# a_1519_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X2 a_1261_n200# a_1061_n264# a_1003_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_n29_n200# a_n229_n264# a_n287_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_229_n200# a_29_n264# a_n29_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_n1319_n200# a_n1519_n264# a_n1577_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_n545_n200# a_n745_n264# a_n803_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_n803_n200# a_n1003_n264# a_n1061_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_n287_n200# a_n487_n264# a_n545_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_n1577_n200# a_n1777_n264# a_n1835_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X10 a_1519_n200# a_1319_n264# a_1261_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_n1061_n200# a_n1261_n264# a_n1319_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X12 a_745_n200# a_545_n264# a_487_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X13 a_1003_n200# a_803_n264# a_745_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_XW23Q2 a_29_n964# a_n2351_n900# a_229_n900# a_n745_n964#
+ a_n1577_n900# a_2035_n900# a_803_n964# a_n2035_n964# a_n545_n900# a_1835_n964# a_1003_n900#
+ a_n229_n964# a_n1003_n964# a_287_n964# a_n2867_n900# a_2093_n964# a_487_n900# a_n29_n900#
+ a_2293_n900# a_1319_n964# a_n1835_n900# a_1061_n964# a_n2293_n964# a_n803_n900#
+ a_1519_n900# a_n2093_n900# a_n1519_n964# a_1261_n900# a_n487_n964# a_n1261_n964#
+ a_2609_n964# a_n1319_n900# a_545_n964# a_n287_n900# a_2351_n964# a_n1061_n900# a_1577_n964#
+ a_2809_n900# a_745_n900# a_n2809_n964# a_2551_n900# a_n2551_n964# w_n3067_n1197#
+ a_1777_n900# a_n2609_n900# a_n1777_n964#
X0 a_1261_n900# a_1061_n964# a_1003_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1 a_n1835_n900# a_n2035_n964# a_n2093_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X2 a_2809_n900# a_2609_n964# a_2551_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X3 a_n2351_n900# a_n2551_n964# a_n2609_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X4 a_n2093_n900# a_n2293_n964# a_n2351_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X5 a_n29_n900# a_n229_n964# a_n287_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X6 a_229_n900# a_29_n964# a_n29_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X7 a_2551_n900# a_2351_n964# a_2293_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X8 a_n1319_n900# a_n1519_n964# a_n1577_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X9 a_n545_n900# a_n745_n964# a_n803_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X10 a_2293_n900# a_2093_n964# a_2035_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X11 a_n803_n900# a_n1003_n964# a_n1061_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X12 a_n287_n900# a_n487_n964# a_n545_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X13 a_n1577_n900# a_n1777_n964# a_n1835_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X14 a_1519_n900# a_1319_n964# a_1261_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X15 a_n1061_n900# a_n1261_n964# a_n1319_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X16 a_745_n900# a_545_n964# a_487_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X17 a_1003_n900# a_803_n964# a_745_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X18 a_487_n900# a_287_n964# a_229_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X19 a_2035_n900# a_1835_n964# a_1777_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X20 a_n2609_n900# a_n2809_n964# a_n2867_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X21 a_1777_n900# a_1577_n964# a_1519_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_RMXH5H a_803_n255# a_1261_n200# a_n1319_n200#
+ a_n287_n200# a_n229_n255# a_n1061_n200# a_287_n255# a_n1003_n255# a_745_n200# a_1319_n255#
+ a_n1711_n422# a_1061_n255# a_229_n200# a_n1577_n200# a_n1519_n255# a_n487_n255#
+ a_n545_n200# a_n1261_n255# a_545_n255# a_1003_n200# a_487_n200# a_n29_n200# a_29_n255#
+ a_n745_n255# a_n803_n200# a_1519_n200#
X0 a_1261_n200# a_1061_n255# a_1003_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_n29_n200# a_n229_n255# a_n287_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_229_n200# a_29_n255# a_n29_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_n1319_n200# a_n1519_n255# a_n1577_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X4 a_n545_n200# a_n745_n255# a_n803_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_n803_n200# a_n1003_n255# a_n1061_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_n287_n200# a_n487_n255# a_n545_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_1519_n200# a_1319_n255# a_1261_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X8 a_n1061_n200# a_n1261_n255# a_n1319_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_745_n200# a_545_n255# a_487_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_1003_n200# a_803_n255# a_745_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_487_n200# a_287_n255# a_229_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NMXZ6U a_n1861_n200# a_n1803_n255# a_n3369_n422#
+ a_n2777_n200# a_n1345_n255# a_n2719_n255# a_2261_n200# a_n1403_n200# a_3177_n200#
+ a_n2319_n200# a_1861_n255# a_2777_n255# a_1403_n255# a_n887_n255# a_n945_n200# a_945_n255#
+ a_2319_n255# a_n487_n200# a_n429_n255# a_1803_n200# a_487_n255# a_2719_n200# a_1345_n200#
+ a_n29_n200# a_n2261_n255# a_887_n200# a_29_n255# a_n3177_n255# a_n3235_n200# a_429_n200#
X0 a_n2319_n200# a_n2719_n255# a_n2777_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X1 a_n2777_n200# a_n3177_n255# a_n3235_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=2
X2 a_2261_n200# a_1861_n255# a_1803_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X3 a_n945_n200# a_n1345_n255# a_n1403_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X4 a_429_n200# a_29_n255# a_n29_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X5 a_1803_n200# a_1403_n255# a_1345_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X6 a_887_n200# a_487_n255# a_429_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X7 a_3177_n200# a_2777_n255# a_2719_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=2
X8 a_n487_n200# a_n887_n255# a_n945_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X9 a_n1403_n200# a_n1803_n255# a_n1861_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X10 a_2719_n200# a_2319_n255# a_2261_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X11 a_n1861_n200# a_n2261_n255# a_n2319_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X12 a_n29_n200# a_n429_n255# a_n487_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X13 a_1345_n200# a_945_n255# a_887_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_BH2H9S a_n229_n1664# a_1061_n1664# a_n1835_n1600#
+ a_n2351_n1600# a_n1261_n1664# a_n1061_n1600# a_1319_n1664# a_1261_n1600# a_287_n1664#
+ a_n2035_n1664# a_2035_n1600# a_n1319_n1600# a_n1519_n1664# a_1519_n1600# a_487_n1600#
+ a_545_n1664# a_29_n1664# a_n487_n1664# a_n287_n1600# w_n2551_n1897# a_745_n1600#
+ a_2093_n1664# a_1577_n1664# a_803_n1664# a_n745_n1664# a_n1003_n1664# a_1003_n1600#
+ a_n545_n1600# a_n2293_n1664# a_n2093_n1600# a_n1777_n1664# a_2293_n1600# a_n1577_n1600#
+ a_1777_n1600# a_n29_n1600# a_1835_n1664# a_229_n1600# a_n803_n1600#
X0 a_n287_n1600# a_n487_n1664# a_n545_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X1 a_n1577_n1600# a_n1777_n1664# a_n1835_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X2 a_n29_n1600# a_n229_n1664# a_n287_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X3 a_2035_n1600# a_1835_n1664# a_1777_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X4 a_n1319_n1600# a_n1519_n1664# a_n1577_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X5 a_n2093_n1600# a_n2293_n1664# a_n2351_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=4.64 ps=32.58 w=16 l=1
X6 a_745_n1600# a_545_n1664# a_487_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X7 a_n1835_n1600# a_n2035_n1664# a_n2093_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X8 a_1261_n1600# a_1061_n1664# a_1003_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X9 a_n545_n1600# a_n745_n1664# a_n803_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X10 a_229_n1600# a_29_n1664# a_n29_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X11 a_1003_n1600# a_803_n1664# a_745_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X12 a_n1061_n1600# a_n1261_n1664# a_n1319_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X13 a_n803_n1600# a_n1003_n1664# a_n1061_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X14 a_1777_n1600# a_1577_n1664# a_1519_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X15 a_1519_n1600# a_1319_n1664# a_1261_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X16 a_487_n1600# a_287_n1664# a_229_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X17 a_2293_n1600# a_2093_n1664# a_2035_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.58 as=2.32 ps=16.29 w=16 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_TT9EEV a_n932_n420# a_1648_n420# a_n1648_n484#
+ a_1390_n420# a_n1390_n484# a_n616_n484# a_n1448_n420# a_674_n484# a_n1190_n420#
+ w_n1906_n717# a_n416_n420# a_874_n420# a_158_n484# a_358_n420# a_n874_n484# a_n1706_n420#
+ a_932_n484# a_100_n420# a_n674_n420# a_1132_n420# a_n358_n484# a_n1132_n484# a_416_n484#
+ a_n158_n420# a_n100_n484# a_616_n420# a_1448_n484# a_1190_n484#
X0 a_n416_n420# a_n616_n484# a_n674_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X1 a_n158_n420# a_n358_n484# a_n416_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X2 a_n1448_n420# a_n1648_n484# a_n1706_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=1.218 ps=8.98 w=4.2 l=1
X3 a_n1190_n420# a_n1390_n484# a_n1448_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X4 a_n674_n420# a_n874_n484# a_n932_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X5 a_n932_n420# a_n1132_n484# a_n1190_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X6 a_358_n420# a_158_n484# a_100_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X7 a_616_n420# a_416_n484# a_358_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X8 a_1648_n420# a_1448_n484# a_1390_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=1.218 pd=8.98 as=0.609 ps=4.49 w=4.2 l=1
X9 a_1132_n420# a_932_n484# a_874_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X10 a_874_n420# a_674_n484# a_616_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X11 a_1390_n420# a_1190_n484# a_1132_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X12 a_100_n420# a_n100_n484# a_n158_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
.ends

.subckt sky130_fd_pr__res_high_po_0p69_XTGLEU a_282_n556# a_282_124# a_516_n556# a_48_124#
+ a_n186_124# a_n420_n556# a_n654_n556# a_516_124# a_48_n556# a_n784_n686# a_n420_124#
+ a_n654_124# a_n186_n556#
X0 a_n420_124# a_n420_n556# a_n784_n686# sky130_fd_pr__res_high_po_0p69 l=1.4
X1 a_48_124# a_48_n556# a_n784_n686# sky130_fd_pr__res_high_po_0p69 l=1.4
X2 a_282_124# a_282_n556# a_n784_n686# sky130_fd_pr__res_high_po_0p69 l=1.4
X3 a_516_124# a_516_n556# a_n784_n686# sky130_fd_pr__res_high_po_0p69 l=1.4
X4 a_n186_124# a_n186_n556# a_n784_n686# sky130_fd_pr__res_high_po_0p69 l=1.4
X5 a_n654_124# a_n654_n556# a_n784_n686# sky130_fd_pr__res_high_po_0p69 l=1.4
.ends

.subckt sky130_td_ip__opamp_hp_narrow avdd vout ibias vinn vinp avss dvdd dvss ena
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_15 avdd avdd m1_n3750_n668# net21 sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_W75H7K_0 net4 avdd net5 net5 avdd net4 avdd net5 net5
+ net5 net5 net3 net5 net5 net3 net4 avdd avdd net5 net5 avdd net4 net3 avdd net5
+ net5 net5 avdd net3 net4 net5 avdd avdd net5 net5 avdd net3 net5 avdd net5 net5
+ net4 net5 net5 avdd net5 net3 avdd net5 net4 avdd net5 net5 avdd net4 net5 net5
+ net5 net4 net5 avdd net3 avdd net5 net3 net5 net4 avdd net3 avdd avdd net5 net5
+ net5 avdd net5 net5 avdd sky130_fd_pr__pfet_g5v0d10v5_W75H7K
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_16 net5 avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_17 m1_n3750_n668# avdd net35 avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_WKXP7K_0 net3 m1_n592_3104# avdd vb2 vb2 net4 m1_n592_3104#
+ vb2 vb2 vb2 vb2 net3 vb2 vb2 net4 net4 net5 net5 vb2 vb2 m1_n592_3104# net3 net3
+ net5 vb2 vb2 vb2 m1_n592_3104# avdd net3 vb2 m1_n592_3104# net5 vb2 vb2 m1_n592_3104#
+ net3 avdd m1_n592_3104# vb2 vb2 net4 vb2 vb2 net5 vb2 avdd avdd avdd net4 net5 vb2
+ net4 net5 vb2 vb2 m1_n592_3104# net3 vb2 vb2 vb2 net3 vb2 m1_n592_3104# net3 m1_n592_3104#
+ vb2 net4 vb2 net4 net5 net4 net5 vb2 vb2 avdd vb2 net5 vb2 avdd vb2 vb2 sky130_fd_pr__pfet_g5v0d10v5_WKXP7K
Xsky130_fd_pr__cap_mim_m3_1_AALY9X_0 net8 m1_n592_3104# m1_32750_1661# m1_n592_3104#
+ net8 m1_32750_1661# m1_32495_1140# m1_32495_1140# m1_n592_3104# net8 m1_32750_1661#
+ m1_32495_1140# sky130_fd_pr__cap_mim_m3_1_AALY9X
Xsky130_fd_pr__nfet_01v8_6H2JYD_0 dvss m1_n6583_10102# m1_n5758_10095# dvss sky130_fd_pr__nfet_01v8_6H2JYD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_0 ibias avss net33 m1_n3750_n668# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_01v8_6H2JYD_1 dvss ena m1_n6583_10102# dvss sky130_fd_pr__nfet_01v8_6H2JYD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_1 net34 avss net31 m1_n3750_n668# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_HQ4STX_0 avdd vb2 vb2 avdd sky130_fd_pr__pfet_g5v0d10v5_HQ4STX
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_2 m1_n3750_n668# avss avss net35 sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_3 net6 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_UKVZ7J_0 net29 avss net12 m1_n4692_n1074# avss m1_n4692_n1074#
+ m1_n4692_n1074# m1_n4692_n1074# avss avss net12 m1_n4692_n1074# m1_n4692_n1074#
+ avss m1_n4692_n1074# m1_n4692_n1074# avss avss net12 avss m1_n4692_n1074# net12
+ avss net12 m1_n4692_n1074# m1_n4692_n1074# avss m1_n4692_n1074# m1_n4692_n1074#
+ avss net29 avss net12 m1_n4692_n1074# net28 m1_n4692_n1074# m1_n4692_n1074# avss
+ net12 m1_n4692_n1074# avss m1_n4692_n1074# avss m1_n4692_n1074# m1_n4692_n1074#
+ net12 m1_n4692_n1074# net28 m1_n4692_n1074# avss avss net12 m1_n4692_n1074# m1_n4692_n1074#
+ sky130_fd_pr__nfet_g5v0d10v5_UKVZ7J
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_4 net10 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_USXRNR_0 avss net10 avss avss avss net6 net5 net10 net10
+ net10 net8 net5 avss net8 net10 net6 avss net10 m1_n592_3104# net6 net10 net6 net5
+ net10 m1_n592_3104# avss net10 avss sky130_fd_pr__nfet_g5v0d10v5_USXRNR
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_0 avdd avdd m1_n3750_n668# net3 sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_5 vb3 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_1 net18 avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_6 m1_n4692_n1074# avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_2 avdd avdd m1_n3750_n668# vb1 sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_7 net33 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_AUMBFF_0 m1_n592_3104# m1_n592_3104# avdd vout avdd
+ vout avdd m1_n592_3104# m1_n592_3104# m1_n592_3104# vout m1_n592_3104# m1_n592_3104#
+ m1_n592_3104# m1_n592_3104# vout m1_n592_3104# m1_n592_3104# m1_n592_3104# avdd
+ avdd avdd avdd m1_n592_3104# m1_n592_3104# avdd vout avdd vout m1_n592_3104# m1_n592_3104#
+ vout avdd m1_n592_3104# vout avdd avdd avdd m1_n592_3104# avdd avdd m1_n592_3104#
+ vout vout m1_n592_3104# m1_n592_3104# vout avdd m1_n592_3104# m1_n592_3104# avdd
+ m1_n592_3104# m1_n592_3104# vout m1_n592_3104# avdd vout avdd m1_n592_3104# m1_n592_3104#
+ vout avdd m1_n592_3104# avdd m1_n592_3104# m1_n592_3104# m1_n592_3104# vout avdd
+ vout sky130_fd_pr__pfet_g5v0d10v5_AUMBFF
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_3 vb5 avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__diode_pw2nd_05v5_25PWK4_0 dvss ena sky130_fd_pr__diode_pw2nd_05v5_25PWK4
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_8 net20 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_4 net13 avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_QL2RRT_0 vinn vinn net1 vinp net1 vtailp vinp vtailp
+ vinp vinn vtailp avdd vinn vtailp vinn avdd vinn vinp net2 avdd vinn avdd vtailp
+ vtailp vinp net1 vtailp vinn net1 vinp net2 vtailp vtailp vinp net2 vinn vinp vinp
+ vinp net2 net1 vtailp vinn net2 vinn net2 avdd vinp vtailp vinn vtailp net1 vtailp
+ vinp sky130_fd_pr__pfet_g5v0d10v5_QL2RRT
Xsky130_fd_pr__cap_mim_m3_2_AALY9W_0 m1_32750_1661# m1_32495_1140# m1_n592_3104# m1_n592_3104#
+ m1_32495_1140# net8 net8 net8 m1_32750_1661# m1_n592_3104# m1_32495_1140# m1_32750_1661#
+ sky130_fd_pr__cap_mim_m3_2_AALY9W
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_9 net31 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_5 avdd avdd m1_n3667_4379# enab_avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_QL2RRT_1 vinp vinp net2 vinn net2 vtailp vinn vtailp
+ vinn vinp vtailp avdd vinp vtailp vinp avdd vinp vinn net1 avdd vinp avdd vtailp
+ vtailp vinn net2 vtailp vinp net2 vinn net1 vtailp vtailp vinn net1 vinp vinn vinn
+ vinn net1 net2 vtailp vinp net1 vinp net1 avdd vinn vtailp vinp vtailp net2 vtailp
+ vinn sky130_fd_pr__pfet_g5v0d10v5_QL2RRT
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_6 avdd avdd m1_n3750_n668# vb2 sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_7 avdd avdd m1_n3750_n668# m1_791_7588# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_01v8_U4BBJH_0 m1_n5758_10095# dvdd m1_n6583_10102# dvdd sky130_fd_pr__pfet_01v8_U4BBJH
Xsky130_fd_pr__pfet_01v8_U4BBJH_1 m1_n6583_10102# dvdd ena dvdd sky130_fd_pr__pfet_01v8_U4BBJH
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_8 m1_180_4838# avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_9 net4 avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_B3XH3Z_0 vtailn avss vb1 avss net12 vb3 vb3 vb3 net29
+ avss vtailn avss net12 vb1 vb3 avss net12 vb3 vb3 net12 net28 avss vtailn vb3 vb3
+ vtailn net12 m1_n4692_n1074# vb3 avss avss vb3 vb3 net12 vb1 vb3 vtailn avss vb3
+ vtailn avss vb3 avss vtailn m1_n4692_n1074# vb3 vb3 net28 vb3 net12 vb3 vb3 vtailn
+ vb3 vtailn vb3 vb3 net12 net29 m1_n4692_n1074# vb3 vb3 sky130_fd_pr__nfet_g5v0d10v5_B3XH3Z
Xsky130_fd_pr__pfet_g5v0d10v5_QTY6KC_0 m1_18668_3467# m1_180_4838# m1_18668_3467#
+ avdd avdd avdd m1_18668_3467# avdd m1_18668_3467# avdd avdd m1_180_4838# m1_180_4838#
+ m1_18668_3467# m1_18668_3467# m1_18668_3467# m1_180_4838# avdd avdd m1_180_4838#
+ avdd avdd m1_18668_3467# m1_180_4838# m1_18668_3467# avdd sky130_fd_pr__pfet_g5v0d10v5_QTY6KC
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_10 net12 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_2B7385_0 avss avss m1_n5910_1250# avss m1_n5910_1250#
+ m1_n5910_1250# m1_n5910_1250# m1_n5910_1250# avss avss m1_n5910_1250# avss avss
+ avss m1_n5910_1250# avss vtailn vtailn m1_n5910_1250# m1_n5910_1250# m1_n5910_1250#
+ vtailn m1_n5910_1250# m1_n5910_1250# m1_n5910_1250# avss vtailn vtailn avss m1_n5910_1250#
+ m1_n5910_1250# avss m1_n5910_1250# avss vtailn vtailn m1_n5910_1250# m1_n5910_1250#
+ sky130_fd_pr__nfet_g5v0d10v5_2B7385
Xsky130_fd_pr__nfet_g5v0d10v5_79TVLH_0 vtailn net4 vtailn vinn vinp net4 net4 vtailn
+ vinn vtailn vinp vtailn vinn vinn vinn avss vinp vtailn vinp net3 vinn avss vinp
+ vtailn vtailn vinn vinp vinp net4 net4 vtailn vinn vinn vtailn net3 vtailn vinn
+ vinp net3 net3 avss vinp net4 vinp vtailn vinp vinn net3 net3 vinp avss avss vtailn
+ vinn sky130_fd_pr__nfet_g5v0d10v5_79TVLH
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_11 net2 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_U73S5M_0 vout vout net8 net8 net8 avss avss vout avss
+ net8 net8 avss vout vout avss net8 net8 net8 net8 net8 net8 avss avss net8 vout
+ avss net8 vout vout avss net8 net8 avss net8 avss avss vout vout net8 avss net8
+ net8 vout net8 net8 net8 net8 net8 net8 net8 avss vout net8 avss avss net8 net8
+ net8 avss vout vout net8 avss net8 vout avss avss vout avss avss sky130_fd_pr__nfet_g5v0d10v5_U73S5M
Xsky130_fd_pr__pfet_g5v0d10v5_PP2RNK_0 vb2 vb1 vtailp avdd vb2 avdd m1_791_7588# vb2
+ vb2 m1_791_7588# avdd vb2 m1_791_7588# vb2 vb2 vb2 vb1 vb2 m1_791_7588# m1_791_7588#
+ vtailp avdd vb2 vb1 vb2 vb2 vtailp m1_791_7588# m1_3549_9621# avdd vtailp vb2 vb2
+ vb2 vtailp vb2 vtailp vb2 m1_791_7588# vb2 vtailp vtailp vb2 m1_791_7588# vb2 avdd
+ vtailp m1_3549_9621# avdd avdd sky130_fd_pr__pfet_g5v0d10v5_PP2RNK
Xsky130_fd_pr__pfet_g5v0d10v5_QTY6H6_0 avdd net22 net22 avdd net22 avdd m1_n3445_8429#
+ avdd net22 avdd net22 avdd net22 m1_n3445_8429# m1_n3445_8429# net22 net22 net22
+ m1_n3445_8429# net32 avdd net22 avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5_QTY6H6
Xsky130_fd_pr__nfet_g5v0d10v5_79TVLH_1 vtailn net3 vtailn vinp vinn net3 net3 vtailn
+ vinp vtailn vinn vtailn vinp vinp vinp avss vinn vtailn vinn net4 vinp avss vinn
+ vtailn vtailn vinp vinn vinn net3 net3 vtailn vinp vinp vtailn net4 vtailn vinp
+ vinn net4 net4 avss vinn net3 vinn vtailn vinn vinp net4 net4 vinn avss avss vtailn
+ vinp sky130_fd_pr__nfet_g5v0d10v5_79TVLH
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_12 net1 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_NT3TPY_0 m1_n5758_10095# net35 avss avss avss avss net35
+ avss avss m1_n3667_4379# m1_n6583_10102# avss m1_n6583_10102# m1_n5758_10095# sky130_fd_pr__nfet_g5v0d10v5_NT3TPY
Xsky130_fd_pr__nfet_g5v0d10v5_5X2ZTR_0 vb2 vb7 vb7 vb7 avss net16 avss vb6 net24 vb7
+ avss vb7 avss net16 vb7 vb6 avss vb7 avss net25 net16 net24 avss vb7 vb6 vb6 vb7
+ vb7 net25 net16 vb2 vb7 vb7 avss net24 net16 vb7 vb2 vb8 vb7 vb7 avss net25 avss
+ vb7 m1_180_4838# net24 avss avss net25 vb7 vb7 vb7 vb2 vb7 m1_180_4838# avss avss
+ vb7 vb7 net25 net24 vb7 vb7 vb7 m1_180_4838# m1_180_4838# vb7 net25 vb7 vb7 vb7
+ net24 vb2 vb7 vb7 vb7 vb7 net16 vb7 vb6 m1_180_4838# sky130_fd_pr__nfet_g5v0d10v5_5X2ZTR
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_13 vb7 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_WK95DB_0 avss net18 vb3 vb3 vb3 vtailn vtailn vb3 vb3
+ net18 net18 vb3 vb3 vtailn vb3 avss net18 avss avss avss net18 vtailn sky130_fd_pr__nfet_g5v0d10v5_WK95DB
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_14 vinp avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_15 m1_n5910_1250# avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_16 vb8 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_PGZBW9_0 net6 net6 net1 net1 avss net6 avss net6 net6
+ avss net6 net6 net6 avss avss net6 net2 net6 avss net6 avss avss net6 net6 net1
+ avss net6 net1 net6 net6 net2 avss avss net6 net6 net2 avss net2 net6 net1 avss
+ net6 net6 net6 net2 net6 net2 avss avss avss avss net1 avss net6 sky130_fd_pr__nfet_g5v0d10v5_PGZBW9
Xsky130_fd_pr__pfet_g5v0d10v5_3QL9S5_0 enab_avdd m1_12266_11884# avdd net21 sky130_fd_pr__pfet_g5v0d10v5_3QL9S5
Xsky130_fd_pr__pfet_g5v0d10v5_U4Z9ZD_1 avdd net35 avdd net35 avdd net35 avdd avdd
+ avdd net35 m1_n3667_4379# avdd avdd avdd m1_n3667_4379# m1_n3667_4379# m1_n3667_4379#
+ m1_n3667_4379# m1_n3667_4379# net35 avdd net35 sky130_fd_pr__pfet_g5v0d10v5_U4Z9ZD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_17 net16 avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_3QL9S5_1 enab_avdd net22 avdd net32 sky130_fd_pr__pfet_g5v0d10v5_3QL9S5
Xsky130_fd_pr__pfet_g5v0d10v5_QSKB8C_0 vb6 vb6 avdd vb3 vb6 vb5 vb6 m1_n4692_n1074#
+ m1_n4692_n1074# vb6 vb6 net13 m1_25484_9858# vb3 vb6 avdd vb6 net10 m1_25484_9858#
+ vb6 vb6 m1_n4692_n1074# vb6 vb6 net13 vb6 vb6 avdd m1_25484_9858# avdd avdd vb6
+ m1_25484_9858# m1_23420_9858# vb6 vb6 m1_n4692_n1074# vb6 vb6 avdd avdd vb6 avdd
+ m1_23420_9858# avdd net10 vb6 vb6 avdd vb6 net13 m1_n4692_n1074# avdd vb6 vb6 vb6
+ avdd m1_25484_9858# vb6 vb6 m1_25484_9858# m1_n4692_n1074# vb3 avdd net10 avdd vb6
+ vb5 vb6 vb5 m1_n4692_n1074# m1_23420_9858# vb6 vb6 vb6 net10 vb3 vb6 sky130_fd_pr__pfet_g5v0d10v5_QSKB8C
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_18 vinn avss avss enab_avdd sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_QRKB8C_0 vb5 vb5 avdd m1_23420_9858# vb5 avdd avdd vb5
+ vb5 avdd vb5 avdd avdd net13 vb5 vb5 avdd m1_25484_9858# avdd avdd avdd m1_25484_9858#
+ vb5 avdd avdd vb5 vb5 avdd vb5 vb5 m1_23420_9858# avdd avdd avdd m1_23420_9858#
+ m1_25484_9858# vb5 vb5 avdd vb5 avdd avdd vb5 net13 vb5 vb5 net13 avdd net13 vb5
+ vb5 vb5 vb5 avdd vb5 vb5 avdd m1_25484_9858# avdd vb5 m1_25484_9858# vb5 vb5 avdd
+ vb5 avdd vb5 avdd avdd vb5 vb5 m1_25484_9858# m1_23420_9858# vb5 sky130_fd_pr__pfet_g5v0d10v5_QRKB8C
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_19 avss avss enab_avdd m1_n3667_4379# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_EVM3FM_0 vb2 vb2 vb2 m1_n5910_1250# vb2 vb2 vtailp vb2
+ avdd vb2 vtailp vb2 avdd m1_n5910_1250# avdd avdd vtailp m1_n5910_1250# m1_n5910_1250#
+ avdd vtailp vtailp sky130_fd_pr__pfet_g5v0d10v5_EVM3FM
Xsky130_fd_pr__nfet_g5v0d10v5_DL2ZHN_0 net16 vb8 vb8 vb8 avss vb8 net24 avss avss
+ vb8 vb8 avss vb8 net25 net16 vb8 vb8 avss avss avss vb8 vb8 net16 net24 vb8 vb8
+ avss avss net16 vb8 vb8 avss avss vb8 net25 net25 vb8 vb8 avss net16 vb8 net24 avss
+ vb8 avss avss vb8 vb8 net24 vb8 net16 vb8 net25 avss vb8 avss avss avss vb8 vb8
+ net24 vb8 avss avss vb8 vb8 avss avss net24 avss vb8 vb8 vb8 avss avss net25 net25
+ avss sky130_fd_pr__nfet_g5v0d10v5_DL2ZHN
Xsky130_fd_pr__nfet_g5v0d10v5_HG2LSW_0 vb3 vb3 avss avss sky130_fd_pr__nfet_g5v0d10v5_HG2LSW
Xsky130_fd_pr__nfet_g5v0d10v5_N64HU4_0 avss avss avss avss ibias net33 net33 avss
+ net20 net20 net20 net34 net33 net33 net33 net33 net21 net33 net33 net20 net33 net21
+ net33 net21 net20 net21 avss avss avss net21 net33 net33 net34 net20 sky130_fd_pr__nfet_g5v0d10v5_N64HU4
Xsky130_fd_pr__nfet_g5v0d10v5_UGZTXE_0 vb3 vb3 net6 net8 net1 avss vb3 net2 vb3 vb3
+ net1 vb3 vb3 vb3 avss net2 avss vb3 net6 vb3 net8 vb3 avss net2 vb3 vb3 net8 net1
+ avss net6 vb3 vb3 net6 net2 net1 vb3 vb3 avss net8 vb3 avss net6 vb3 net6 net1 avss
+ vb3 vb3 net8 vb3 net8 net6 vb3 net2 net2 net8 net1 vb3 sky130_fd_pr__nfet_g5v0d10v5_UGZTXE
Xsky130_fd_pr__pfet_g5v0d10v5_Q46EE6_0 m1_n3445_8429# m1_12266_11884# m1_12266_11884#
+ avdd net21 m1_12266_11884# m1_n3445_8429# net32 avdd m1_n3445_8429# avdd avdd m1_12266_11884#
+ m1_n3445_8429# avdd net32 m1_12266_11884# vb7 vb7 m1_12266_11884# avdd m1_12266_11884#
+ vb7 vb7 m1_12266_11884# avdd m1_12266_11884# avdd vb7 m1_12266_11884# sky130_fd_pr__pfet_g5v0d10v5_Q46EE6
Xsky130_fd_pr__pfet_g5v0d10v5_XW23Q2_0 vb1 m1_791_7588# m1_3549_9621# vb1 avdd avdd
+ vb1 vb1 avdd vb1 avdd vb1 vb1 vb1 avdd vb1 avdd avdd m1_791_7588# vb1 m1_791_7588#
+ vb1 vb1 m1_791_7588# avdd avdd vb1 m1_791_7588# vb1 vb1 avdd m1_791_7588# vb1 m1_3549_9621#
+ vb1 avdd vb1 avdd m1_791_7588# avdd avdd vb1 avdd m1_791_7588# avdd vb1 sky130_fd_pr__pfet_g5v0d10v5_XW23Q2
Xsky130_fd_pr__nfet_g5v0d10v5_RMXH5H_0 m1_18790_1436# avss net10 net10 avss m1_18790_1436#
+ m1_18790_1436# net10 avss avss avss m1_18790_1436# avss avss avss net10 m1_18790_1436#
+ net10 m1_18790_1436# m1_18790_1436# m1_18790_1436# avss avss net10 net10 avss sky130_fd_pr__nfet_g5v0d10v5_RMXH5H
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_10 net32 avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_NMXZ6U_0 net20 net31 avss net20 net31 net31 avss avss
+ avss avss net31 avss net31 net31 net20 net31 net31 avss net31 net20 net31 net20
+ avss net34 net31 net20 net31 avss avss avss sky130_fd_pr__nfet_g5v0d10v5_NMXZ6U
Xsky130_fd_pr__pfet_g5v0d10v5_BH2H9S_0 net18 net18 vtailp avdd net18 avdd net18 vtailp
+ net18 net18 avdd vtailp net18 avdd avdd net18 net18 net18 net18 avdd vtailp avdd
+ net18 net18 net18 net18 avdd avdd avdd avdd net18 avdd avdd vtailp avdd net18 net18
+ vtailp sky130_fd_pr__pfet_g5v0d10v5_BH2H9S
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_11 net22 avdd m1_n3750_n668# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_TT9EEV_0 net5 avdd avdd net8 m1_180_4838# m1_180_4838#
+ net5 m1_180_4838# net6 avdd net5 net8 avdd avdd m1_180_4838# avdd m1_180_4838# net5
+ net6 m1_n592_3104# m1_180_4838# m1_180_4838# avdd net6 m1_180_4838# m1_n592_3104#
+ avdd m1_180_4838# sky130_fd_pr__pfet_g5v0d10v5_TT9EEV
Xsky130_fd_pr__res_high_po_0p69_XTGLEU_0 m1_32032_n77# m1_32750_1661# avss m1_32495_1140#
+ vout m1_32032_n77# avss avss m1_32268_124# avss vout avss m1_32268_124# sky130_fd_pr__res_high_po_0p69_XTGLEU
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_12 avdd avdd m1_n3750_n668# vb6 sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13 avdd avdd m1_n3750_n668# m1_n592_3104# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_14 avdd avdd m1_n3750_n668# m1_n3445_8429# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
.ends

.subckt sky130_fd_sc_hvl__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.4275 ps=3.57 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.21375 ps=2.07 w=0.75 l=0.5
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP a_214_n1416# a_n118_984# a_48_n1416#
+ a_n450_984# a_n580_n1546# a_n284_n1416# a_n118_n1416# a_48_984# a_380_984# a_380_n1416#
+ a_214_984# a_n284_984# a_n450_n1416#
X0 a_n118_984# a_n118_n1416# a_n580_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X1 a_380_984# a_380_n1416# a_n580_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X2 a_214_984# a_214_n1416# a_n580_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X3 a_n284_984# a_n284_n1416# a_n580_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X4 a_n450_984# a_n450_n1416# a_n580_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X5 a_48_984# a_48_n1416# a_n580_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_92HZNS a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_TUFYNQ a_n50_n197# a_50_n100# w_n308_n397# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n308_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt T_Gate_5V UPPER PGATE NGATE LOWER AVSS AVDD
XXM1 LOWER AVSS UPPER NGATE sky130_fd_pr__nfet_g5v0d10v5_92HZNS
XXM2 PGATE LOWER AVDD UPPER sky130_fd_pr__pfet_g5v0d10v5_TUFYNQ
.ends

.subckt Universal_R_2R_Block2 VD DVDD VIRTOUT CMOUT R2RIN R2ROUT AVSS DVSS AVDD
Xx1 VD DVDD DVSS AVDD AVDD VDbuf AVDD DVSS DVSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xx2 VDbuf DVSS DVSS AVDD AVDD VDBAR sky130_fd_sc_hvl__inv_1
Xsky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_0 m1_4390_n2466# m1_6792_n1970# m1_4394_n2136#
+ x13/LOWER AVSS m1_4392_n1802# m1_4394_n2136# R2ROUT R2RIN m1_4390_n2466# R2ROUT
+ m1_6792_n1970# m1_4392_n1802# sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP
Xsky130_fd_sc_hvl__diode_2_0 VD DVSS DVSS AVDD AVDD sky130_fd_sc_hvl__diode_2
Xx12 VIRTOUT VDBAR VDbuf x13/LOWER AVSS AVDD T_Gate_5V
Xx13 CMOUT VDbuf VDBAR x13/LOWER AVSS AVDD T_Gate_5V
.ends

.subckt sky130_fd_pr__res_high_po_0p69_FJD3D2 a_n199_n4646# a_n69_4084# a_n69_n4516#
X0 a_n69_4084# a_n69_n4516# a_n199_n4646# sky130_fd_pr__res_high_po_0p69 l=41
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_FEJX3A a_952_n991# a_n1352_n573# a_200_318# a_318_736#
+ a_n952_n518# a_n258_n100# a_n952_736# a_776_n100# a_n834_318# a_n776_n991# a_n258_n936#
+ a_n258_736# a_952_681# a_776_n936# a_894_736# a_n834_n518# a_n200_n573# a_318_n100#
+ a_776_318# a_200_n518# a_n1352_681# a_376_n991# a_1352_n518# a_318_n936# a_n376_n518#
+ a_894_n518# a_318_318# a_n1544_n1158# a_952_n573# a_n1352_n155# a_n952_318# a_n1410_n100#
+ a_n1410_736# a_n376_736# a_n200_681# a_n1410_n936# a_n258_n518# a_n776_n573# a_n258_318#
+ a_776_n518# a_894_318# a_952_263# a_n200_n155# a_1352_736# a_376_681# a_n1352_263#
+ a_318_n518# a_376_n573# a_n776_681# a_n952_n100# a_952_n155# a_200_736# a_n952_n936#
+ a_n1352_n991# a_n1410_318# a_n376_318# a_n200_263# a_n776_n155# a_n834_736# a_n1410_n518#
+ a_n834_n100# a_200_n100# a_1352_318# a_n200_n991# a_1352_n100# a_376_263# a_n834_n936#
+ a_n376_n100# a_776_736# a_1352_n936# a_200_n936# a_894_n100# a_376_n155# a_n376_n936#
+ a_n776_263# a_894_n936#
X0 a_1352_n518# a_952_n573# a_894_n518# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X1 a_n376_n518# a_n776_n573# a_n834_n518# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X2 a_n952_n100# a_n1352_n155# a_n1410_n100# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X3 a_n376_n100# a_n776_n155# a_n834_n100# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X4 a_200_n100# a_n200_n155# a_n258_n100# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X5 a_776_736# a_376_681# a_318_736# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X6 a_1352_736# a_952_681# a_894_736# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X7 a_n952_n518# a_n1352_n573# a_n1410_n518# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X8 a_n952_318# a_n1352_263# a_n1410_318# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X9 a_776_n936# a_376_n991# a_318_n936# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X10 a_200_n936# a_n200_n991# a_n258_n936# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X11 a_n376_318# a_n776_263# a_n834_318# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X12 a_200_318# a_n200_263# a_n258_318# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X13 a_776_n100# a_376_n155# a_318_n100# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X14 a_1352_n100# a_952_n155# a_894_n100# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X15 a_n376_n936# a_n776_n991# a_n834_n936# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X16 a_1352_n936# a_952_n991# a_894_n936# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X17 a_776_318# a_376_263# a_318_318# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X18 a_1352_318# a_952_263# a_894_318# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X19 a_n952_n936# a_n1352_n991# a_n1410_n936# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X20 a_n952_736# a_n1352_681# a_n1410_736# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X21 a_200_736# a_n200_681# a_n258_736# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X22 a_776_n518# a_376_n573# a_318_n518# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X23 a_n376_736# a_n776_681# a_n834_736# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
X24 a_200_n518# a_n200_n573# a_n258_n518# a_n1544_n1158# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NZU856 a_616_n1610# a_n2938_n2808# a_n2738_n500#
+ a_874_n2720# a_n1190_n1610# a_1132_1720# a_n1448_610# a_n932_610# a_n416_n1610#
+ a_1390_n1610# a_1906_n500# a_n674_n2720# a_1132_n2720# a_n2480_n500# a_n2996_1720#
+ a_n2164_n2808# a_n416_610# a_n2738_n1610# a_n2996_n2720# a_1390_610# a_2938_n1610#
+ a_n1648_n2808# a_358_n500# a_n158_1720# a_2222_n2808# a_2164_n500# a_874_610# a_1706_n2808#
+ a_n1706_n500# a_2164_n1610# a_674_n2808# a_n674_n500# a_100_n500# a_n1448_n1610#
+ a_358_610# a_616_1720# a_1648_n1610# a_n1964_1720# a_2422_1720# a_n100_n2808# a_n932_n2720#
+ a_n1190_610# a_358_n2720# a_n932_1720# a_1132_n500# a_100_n1610# a_n158_n2720# a_n2422_n2808#
+ a_1648_1720# a_n674_610# a_n1906_n2808# a_n2996_n500# a_1390_1720# a_n158_610# a_n2222_1720#
+ a_n2222_n1610# a_n2480_n2720# a_n158_n500# a_2422_n1610# a_2680_n2720# a_932_n2808#
+ a_n1132_n2808# a_n1706_n1610# a_n874_n2808# a_n1964_n2720# a_n1448_1720# a_1906_n1610#
+ a_158_n2808# a_874_n1610# a_616_n2720# a_n1190_1720# a_616_n500# a_n674_n1610# a_n1190_n2720#
+ a_n416_1720# a_2938_610# a_2422_610# a_n1964_n500# a_1132_n1610# a_1390_n2720# a_n416_n2720#
+ a_1906_610# a_2422_n500# a_2938_1720# a_n2996_n1610# a_874_1720# a_n2738_n2720#
+ a_n932_n500# a_2938_n2720# a_2480_n2808# a_2680_1720# a_1648_n500# a_1964_n2808#
+ a_n2222_n500# a_1390_n500# a_n2738_1720# a_2164_n2720# a_416_n2808# a_n358_n2808#
+ a_n2738_610# a_n1448_n2720# a_n2222_610# a_n1706_610# a_1648_n2720# a_1906_1720#
+ a_1190_n2808# a_n2480_1720# a_n1448_n500# a_n932_n1610# a_358_n1610# a_2680_610#
+ a_n2680_n2808# a_n158_n1610# a_358_1720# a_n1190_n500# a_2738_n2808# a_2164_610#
+ a_100_n2720# a_n416_n500# a_1648_610# a_2164_1720# a_1132_610# a_n1706_1720# a_2938_n500#
+ a_874_n500# a_n2480_n1610# a_100_1720# a_n674_1720# a_2680_n1610# a_n2222_n2720#
+ a_n1390_n2808# a_100_610# a_616_610# a_n1964_n1610# a_2680_n500# a_1448_n2808# a_2422_n2720#
+ a_n616_n2808# a_n3130_n2942# a_n1706_n2720# a_n2996_610# a_n2480_610# a_1906_n2720#
+ a_n1964_610#
X0 a_n2480_n2720# a_n2680_n2808# a_n2738_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X1 a_n1448_n1610# a_n1648_n2808# a_n1706_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_2938_n2720# a_2738_n2808# a_2680_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X3 a_1906_n1610# a_1706_n2808# a_1648_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a_1906_n500# a_1706_n2808# a_1648_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X5 a_1648_n500# a_1448_n2808# a_1390_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X6 a_1906_1720# a_1706_n2808# a_1648_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X7 a_n1190_n2720# a_n1390_n2808# a_n1448_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X8 a_1648_1720# a_1448_n2808# a_1390_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X9 a_2938_610# a_2738_n2808# a_2680_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X10 a_n674_610# a_n874_n2808# a_n932_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X11 a_1648_n2720# a_1448_n2808# a_1390_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X12 a_n1448_610# a_n1648_n2808# a_n1706_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X13 a_n1964_610# a_n2164_n2808# a_n2222_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X14 a_874_n1610# a_674_n2808# a_616_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X15 a_2680_n1610# a_2480_n2808# a_2422_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X16 a_1132_n500# a_932_n2808# a_874_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X17 a_1132_1720# a_932_n2808# a_874_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X18 a_n1964_n1610# a_n2164_n2808# a_n2222_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X19 a_874_n500# a_674_n2808# a_616_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X20 a_1390_610# a_1190_n2808# a_1132_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X21 a_616_n1610# a_416_n2808# a_358_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X22 a_874_1720# a_674_n2808# a_616_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X23 a_2422_n1610# a_2222_n2808# a_2164_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X24 a_1390_n1610# a_1190_n2808# a_1132_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X25 a_n2738_610# a_n2938_n2808# a_n2996_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X26 a_358_n2720# a_158_n2808# a_100_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X27 a_n674_n1610# a_n874_n2808# a_n932_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X28 a_2164_610# a_1964_n2808# a_1906_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X29 a_2164_n500# a_1964_n2808# a_1906_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X30 a_2680_610# a_2480_n2808# a_2422_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X31 a_n416_n1610# a_n616_n2808# a_n674_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X32 a_616_610# a_416_n2808# a_358_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X33 a_2164_1720# a_1964_n2808# a_1906_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X34 a_n2738_n500# a_n2938_n2808# a_n2996_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X35 a_100_n2720# a_n100_n2808# a_n158_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X36 a_n2738_n2720# a_n2938_n2808# a_n2996_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X37 a_n1706_n1610# a_n1906_n2808# a_n1964_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X38 a_n2738_1720# a_n2938_n2808# a_n2996_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X39 a_n158_n2720# a_n358_n2808# a_n416_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X40 a_n2480_n500# a_n2680_n2808# a_n2738_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X41 a_n1190_610# a_n1390_n2808# a_n1448_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X42 a_1390_n500# a_1190_n2808# a_1132_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X43 a_n2480_1720# a_n2680_n2808# a_n2738_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X44 a_2164_n2720# a_1964_n2808# a_1906_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X45 a_n2222_n500# a_n2422_n2808# a_n2480_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X46 a_1390_1720# a_1190_n2808# a_1132_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X47 a_n1448_n2720# a_n1648_n2808# a_n1706_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X48 a_n2222_1720# a_n2422_n2808# a_n2480_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X49 a_n1964_n500# a_n2164_n2808# a_n2222_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X50 a_1906_n2720# a_1706_n2808# a_1648_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X51 a_n1964_1720# a_n2164_n2808# a_n2222_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X52 a_1132_n1610# a_932_n2808# a_874_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X53 a_n2480_610# a_n2680_n2808# a_n2738_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X54 a_n2222_n1610# a_n2422_n2808# a_n2480_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X55 a_100_n500# a_n100_n2808# a_n158_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X56 a_874_n2720# a_674_n2808# a_616_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X57 a_100_1720# a_n100_n2808# a_n158_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X58 a_2680_n2720# a_2480_n2808# a_2422_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X59 a_n1964_n2720# a_n2164_n2808# a_n2222_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X60 a_n932_n1610# a_n1132_n2808# a_n1190_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X61 a_358_610# a_158_n2808# a_100_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X62 a_616_n2720# a_416_n2808# a_358_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X63 a_2422_n2720# a_2222_n2808# a_2164_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X64 a_1390_n2720# a_1190_n2808# a_1132_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X65 a_2938_n500# a_2738_n2808# a_2680_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X66 a_1132_610# a_932_n2808# a_874_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X67 a_2938_1720# a_2738_n2808# a_2680_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X68 a_n416_610# a_n616_n2808# a_n674_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X69 a_n674_n2720# a_n874_n2808# a_n932_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X70 a_2422_n500# a_2222_n2808# a_2164_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X71 a_n416_n500# a_n616_n2808# a_n674_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X72 a_2422_1720# a_2222_n2808# a_2164_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X73 a_n416_n2720# a_n616_n2808# a_n674_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X74 a_n158_n500# a_n358_n2808# a_n416_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X75 a_n416_1720# a_n616_n2808# a_n674_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X76 a_n158_1720# a_n358_n2808# a_n416_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X77 a_n1706_n2720# a_n1906_n2808# a_n1964_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X78 a_n2480_n1610# a_n2680_n2808# a_n2738_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X79 a_2938_n1610# a_2738_n2808# a_2680_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X80 a_n1190_n1610# a_n1390_n2808# a_n1448_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X81 a_1906_610# a_1706_n2808# a_1648_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X82 a_1648_n1610# a_1448_n2808# a_1390_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X83 a_2422_610# a_2222_n2808# a_2164_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X84 a_1132_n2720# a_932_n2808# a_874_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X85 a_n932_610# a_n1132_n2808# a_n1190_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X86 a_874_610# a_674_n2808# a_616_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X87 a_n1706_n500# a_n1906_n2808# a_n1964_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X88 a_n158_610# a_n358_n2808# a_n416_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X89 a_n2222_n2720# a_n2422_n2808# a_n2480_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X90 a_2680_n500# a_2480_n2808# a_2422_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X91 a_n1706_1720# a_n1906_n2808# a_n1964_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X92 a_n1448_n500# a_n1648_n2808# a_n1706_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X93 a_n674_n500# a_n874_n2808# a_n932_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X94 a_n1190_n500# a_n1390_n2808# a_n1448_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X95 a_n1448_1720# a_n1648_n2808# a_n1706_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X96 a_2680_1720# a_2480_n2808# a_2422_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X97 a_n674_1720# a_n874_n2808# a_n932_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X98 a_n932_n2720# a_n1132_n2808# a_n1190_n2720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X99 a_n1190_1720# a_n1390_n2808# a_n1448_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X100 a_100_610# a_n100_n2808# a_n158_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X101 a_n1706_610# a_n1906_n2808# a_n1964_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X102 a_358_n1610# a_158_n2808# a_100_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X103 a_n932_n500# a_n1132_n2808# a_n1190_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X104 a_n932_1720# a_n1132_n2808# a_n1190_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X105 a_n2222_610# a_n2422_n2808# a_n2480_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X106 a_616_n500# a_416_n2808# a_358_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X107 a_616_1720# a_416_n2808# a_358_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X108 a_358_n500# a_158_n2808# a_100_n500# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X109 a_100_n1610# a_n100_n2808# a_n158_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X110 a_n2738_n1610# a_n2938_n2808# a_n2996_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X111 a_1648_610# a_1448_n2808# a_1390_610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X112 a_358_1720# a_158_n2808# a_100_1720# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X113 a_n158_n1610# a_n358_n2808# a_n416_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X114 a_2164_n1610# a_1964_n2808# a_1906_n1610# a_n3130_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_AJ3MPE a_72_772# a_n90_n750# a_n138_n838# a_n182_n750#
+ a_n284_n924# a_120_n750# a_28_n750#
X0 a_120_n750# a_72_772# a_28_n750# a_n284_n924# sky130_fd_pr__nfet_01v8_lvt ad=2.325 pd=15.62 as=2.325 ps=15.62 w=7.5 l=0.15
X1 a_n90_n750# a_n138_n838# a_n182_n750# a_n284_n924# sky130_fd_pr__nfet_01v8_lvt ad=2.325 pd=15.62 as=2.325 ps=15.62 w=7.5 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_UX3DP3 a_n1087_n4118# a_29_n4215# a_1029_118#
+ a_n29_n4118# a_29_21# a_n1029_21# w_n1225_n4337# a_n1087_118# a_1029_n4118# a_n1029_n4215#
+ a_n29_118#
X0 a_n29_n4118# a_n1029_n4215# a_n1087_n4118# w_n1225_n4337# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=5.8 ps=40.58 w=20 l=5
X1 a_1029_n4118# a_29_n4215# a_n29_n4118# w_n1225_n4337# sky130_fd_pr__pfet_01v8_lvt ad=5.8 pd=40.58 as=2.9 ps=20.29 w=20 l=5
X2 a_1029_118# a_29_21# a_n29_118# w_n1225_n4337# sky130_fd_pr__pfet_01v8_lvt ad=5.8 pd=40.58 as=2.9 ps=20.29 w=20 l=5
X3 a_n29_118# a_n1029_21# a_n1087_118# w_n1225_n4337# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=5.8 ps=40.58 w=20 l=5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_8UL4MK a_467_n1000# a_n803_n1000# w_n1559_n1297#
+ a_1301_n1000# a_n645_n1000# a_1143_n1000# a_189_n1000# a_n525_n1000# a_923_n1097#
+ a_1023_n1000# a_n1201_n1000# a_n367_n1000# a_n1359_n1000# a_n745_n1097# a_n89_n1000#
+ a_n247_n1000# a_645_n1097# a_865_n1000# a_n467_n1097# a_n1301_n1097# a_745_n1000#
+ a_n1081_n1000# a_367_n1097# a_89_n1097# a_587_n1000# a_309_n1000# a_31_n1000# a_n923_n1000#
+ a_1201_n1097# a_n189_n1097# a_n1023_n1097#
X0 a_n1201_n1000# a_n1301_n1097# a_n1359_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X1 a_1301_n1000# a_1201_n1097# a_1143_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X2 a_189_n1000# a_89_n1097# a_31_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X3 a_n645_n1000# a_n745_n1097# a_n803_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X4 a_745_n1000# a_645_n1097# a_587_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X5 a_n89_n1000# a_n189_n1097# a_n247_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X6 a_n923_n1000# a_n1023_n1097# a_n1081_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X7 a_1023_n1000# a_923_n1097# a_865_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X8 a_n367_n1000# a_n467_n1097# a_n525_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
X9 a_467_n1000# a_367_n1097# a_309_n1000# w_n1559_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.5
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_BHK9HY c1_n3758_n5640# c1_1466_n5640# m3_1426_n5680#
+ m3_n1186_n5680# m3_n3798_n5680# c1_n1146_n5640#
X0 c1_n3758_n5640# m3_n3798_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X1 c1_n1146_n5640# m3_n1186_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X2 c1_1466_n5640# m3_1426_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X3 c1_n3758_n5640# m3_n3798_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X4 c1_1466_n5640# m3_1426_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X5 c1_n3758_n5640# m3_n3798_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X6 c1_n1146_n5640# m3_n1186_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X7 c1_n3758_n5640# m3_n3798_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X8 c1_n1146_n5640# m3_n1186_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X9 c1_1466_n5640# m3_1426_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X10 c1_1466_n5640# m3_1426_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X11 c1_1466_n5640# m3_1426_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X12 c1_n1146_n5640# m3_n1186_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X13 c1_n3758_n5640# m3_n3798_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X14 c1_n1146_n5640# m3_n1186_n5680# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
.ends

.subckt x1_x32_OA VDD VOUT VINN VINP VBIAS w_8718_n902# w_7736_n902# VSS w_4240_n902#
XXR1 VSS m1_10706_1822# VOUT sky130_fd_pr__res_high_po_0p69_FJD3D2
Xsky130_fd_pr__nfet_05v0_nvt_FEJX3A_0 VINP VINP w_8718_n902# w_8718_n902# w_8718_n902#
+ m1_9368_n744# w_8718_n902# m1_9368_n744# w_8718_n902# VINP m1_9368_n744# m1_9368_n744#
+ VINP m1_9368_n744# m1_9368_n744# w_8718_n902# VINP w_8718_n902# m1_9368_n744# w_8718_n902#
+ VINP VINP w_8718_n902# w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902# w_8718_n902#
+ VINP VINP w_8718_n902# m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP m1_9368_n744#
+ m1_9368_n744# VINP m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902#
+ VINP VINP w_8718_n902# VINP VINP w_8718_n902# VINP w_8718_n902# w_8718_n902# VINP
+ m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902# m1_9368_n744# w_8718_n902# w_8718_n902#
+ w_8718_n902# VINP w_8718_n902# VINP w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902#
+ w_8718_n902# m1_9368_n744# VINP m1_9368_n744# VINP m1_9368_n744# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
Xsky130_fd_pr__nfet_g5v0d10v5_NZU856_0 VSS VBIAS VOUT VOUT VOUT VSS VSS VSS VSS VOUT
+ VOUT VOUT VSS VSS VSS VBIAS VSS VOUT VSS VOUT w_7736_n902# VBIAS VOUT VOUT VBIAS
+ VSS VOUT VBIAS VOUT VSS VBIAS VOUT VSS VSS VOUT VSS VSS VSS w_7736_n902# VBIAS VSS
+ VOUT VOUT VSS VSS VSS VOUT VBIAS VSS VOUT VBIAS VSS VOUT VOUT VOUT VOUT VSS VOUT
+ w_7736_n902# VSS VBIAS VBIAS VOUT VBIAS VSS VSS VOUT VBIAS VOUT VSS VOUT VSS VOUT
+ VOUT VSS w_7736_n902# w_7736_n902# VSS VSS VOUT VSS VOUT w_7736_n902# w_7736_n902#
+ VSS VOUT VOUT VSS w_7736_n902# VBIAS VSS VSS VBIAS VOUT VOUT VOUT VSS VBIAS VBIAS
+ VOUT VSS VOUT VOUT VSS VOUT VBIAS VSS VSS VSS VOUT VSS VBIAS VOUT VOUT VOUT VBIAS
+ VSS VSS VSS VSS VSS VSS VOUT w_7736_n902# VOUT VSS VSS VOUT VSS VOUT VBIAS VSS VSS
+ VSS VSS VBIAS w_7736_n902# VBIAS VSS VOUT VSS VSS VOUT VSS sky130_fd_pr__nfet_g5v0d10v5_NZU856
XXM2 VINN w_8718_n902# VINP w_7736_n902# w_7736_n902# w_4240_n902# w_7736_n902# sky130_fd_pr__nfet_01v8_lvt_AJ3MPE
XXM6 m1_9368_n744# m1_4902_n766# m1_9368_n744# VDD m1_4902_n766# m1_4902_n766# VDD
+ m1_4902_n766# m1_4902_n766# m1_4902_n766# VDD sky130_fd_pr__pfet_01v8_lvt_UX3DP3
XXM8 VDD VOUT VDD VOUT VDD VDD VOUT VDD m1_9368_n744# VDD VDD VOUT VOUT m1_9368_n744#
+ VDD VOUT m1_9368_n744# VOUT m1_9368_n744# m1_9368_n744# VOUT VDD m1_9368_n744# m1_9368_n744#
+ VDD VOUT VDD VOUT m1_9368_n744# m1_9368_n744# m1_9368_n744# sky130_fd_pr__pfet_g5v0d10v5_8UL4MK
Xsky130_fd_pr__cap_mim_m3_1_BHK9HY_0 m1_9368_n744# m1_9368_n744# m1_10706_1822# m1_10706_1822#
+ m1_10706_1822# m1_9368_n744# sky130_fd_pr__cap_mim_m3_1_BHK9HY
XXM10 VINN VINN m1_4902_n766# m1_4902_n766# m1_4902_n766# w_4240_n902# m1_4902_n766#
+ w_4240_n902# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902#
+ m1_4902_n766# VINN m1_4902_n766# w_4240_n902# m1_4902_n766# VINN VINN m1_4902_n766#
+ m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# w_4240_n902# VINN VINN m1_4902_n766#
+ w_4240_n902# w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902#
+ w_4240_n902# w_4240_n902# VINN VINN m1_4902_n766# VINN VINN m1_4902_n766# VINN VINN
+ m1_4902_n766# VINN m1_4902_n766# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN
+ VINN m1_4902_n766# w_4240_n902# m1_4902_n766# m1_4902_n766# m1_4902_n766# VINN m1_4902_n766#
+ VINN m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# m1_4902_n766# w_4240_n902#
+ VINN w_4240_n902# VINN w_4240_n902# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_3WU84W a_n3899_n1610# a_n29_n2720# a_3067_1720#
+ a_4357_n2720# a_1261_n500# a_n287_610# a_n4673_610# a_487_n1610# a_1777_1720# a_n2609_1720#
+ a_4873_1720# a_n803_n2720# a_n3641_610# a_n5705_1720# a_n5389_n2808# a_229_n2720#
+ a_3383_n2808# a_n5189_610# a_n287_n1610# a_n3641_n2720# a_n4157_610# a_2867_n2808#
+ a_3841_n2720# a_n2351_1720# a_n1319_n500# a_5389_1720# a_3583_n500# a_n3125_610#
+ a_5447_n2808# a_n4415_n500# a_n5705_n2720# a_n2609_610# a_n4873_n2808# a_3067_n2720#
+ a_n287_n500# a_229_1720# a_n5189_n1610# a_n1061_n500# a_4099_n500# a_3583_610# a_n1577_1720#
+ a_5389_n1610# a_n4099_n2808# a_n4673_1720# a_4931_n2808# a_2093_n2808# a_2551_610#
+ a_2035_1720# a_n2351_n2720# a_4099_610# a_5131_1720# a_1577_n2808# a_2551_n2720#
+ a_803_n2808# a_n745_n2808# a_n1003_n2808# a_n4673_n1610# a_n1835_n2720# a_2809_n500#
+ a_3067_610# a_3841_1720# a_4157_n2808# a_5131_n2720# a_745_n500# a_n5189_1720# a_4873_n1610#
+ a_n4415_n2720# a_n3383_n500# a_2035_610# a_n545_1720# a_n3899_1720# a_n3583_n2808#
+ a_4615_n2720# a_1519_610# a_1003_610# a_745_n1610# a_4357_1720# a_2551_n500# a_4099_n1610#
+ a_3641_n2808# a_n5647_n2808# a_n1061_n2720# a_n545_n1610# a_1003_n1610# a_1261_n2720#
+ a_n3383_n1610# a_3067_n500# a_1777_n500# a_n3899_610# a_n3641_1720# a_3583_n1610#
+ a_n2609_n500# a_n3383_610# a_1003_1720# a_n2293_n2808# a_4873_n500# a_n2867_n1610#
+ a_n3125_n2720# a_n5705_n500# a_n2351_610# a_n2867_610# a_3325_n2720# a_n5447_n1610#
+ a_n2609_n2720# a_n1835_610# a_n1777_n2808# a_5647_n1610# a_n4157_1720# a_n4357_n2808#
+ a_2809_n2720# a_n2351_n500# a_2351_n2808# a_5389_n500# a_n2867_1720# a_n1319_610#
+ a_3325_1720# a_1835_n2808# a_n803_610# a_n4931_n1610# a_n2093_n1610# a_229_n500#
+ a_4415_n2808# a_2293_n1610# a_n3841_n2808# a_n1577_n1610# a_n1577_n500# a_n5705_610#
+ a_n4673_n500# a_2293_610# a_2035_n2720# a_n229_n2808# a_n4157_n1610# a_n29_n1610#
+ a_1777_n1610# a_n1319_n2720# a_2035_n500# a_1777_610# a_1261_610# a_n29_1720# a_5131_n500#
+ a_4357_n1610# a_1519_n2720# a_5647_1720# a_487_1720# a_n3067_n2808# a_3841_n500#
+ a_1061_n2808# a_n3899_n2720# a_n803_n1610# a_n5189_n500# a_229_n1610# a_n545_n500#
+ a_487_n2720# a_n3899_n500# a_n3641_n1610# a_2293_1720# a_n3125_1720# a_745_610#
+ a_3125_n2808# a_4357_n500# a_n1835_1720# a_3841_n1610# a_n4931_1720# a_n2551_n2808#
+ a_n287_n2720# a_5647_610# a_5131_610# a_2609_n2808# a_4615_610# a_n5131_n2808# a_n5705_n1610#
+ a_229_610# a_3067_n1610# a_n4615_n2808# a_n5447_1720# a_n3641_n500# a_n803_1720#
+ a_n5189_n2720# a_1003_n500# a_n2093_610# a_1519_1720# a_n2351_n1610# a_5389_n2720#
+ a_n1577_610# a_4615_1720# a_n1061_610# a_n2093_1720# a_2551_n1610# a_n4157_n500#
+ a_n1261_n2808# a_n1835_n1610# a_1319_n2808# a_5131_n1610# a_n2867_n500# a_n4415_n1610#
+ a_1261_1720# a_n4673_n2720# a_n545_610# a_3325_n500# a_n4931_610# a_3899_n2808#
+ a_4615_n1610# a_4873_n2720# a_287_n2808# a_n3325_n2808# a_n5447_610# a_n2809_n2808#
+ a_745_n2720# a_n1061_n1610# a_4099_n2720# a_n4415_610# a_n1319_1720# a_n29_n500#
+ a_3583_1720# a_n4415_1720# a_1261_n1610# a_5647_n500# a_n545_n2720# a_487_n500#
+ a_1003_n2720# a_n287_1720# a_n3125_n1610# a_n3383_n2720# a_4873_610# a_n1061_1720#
+ a_4099_1720# a_3325_n1610# a_3583_n2720# a_2293_n500# a_n3125_n500# a_487_610# a_n2035_n2808#
+ a_n2609_n1610# a_n2867_n2720# a_3841_610# a_5189_n2808# a_n1835_n500# a_2809_n1610#
+ a_n4931_n500# a_5389_610# a_n1519_n2808# a_n5447_n2720# a_4357_610# a_5647_n2720#
+ a_2809_1720# a_n29_610# a_3325_610# a_745_1720# a_n3383_1720# a_n5447_n500# a_2809_610#
+ a_4673_n2808# a_n5839_n2942# a_n4931_n2720# a_n2093_n2720# a_n803_n500# a_2551_1720#
+ a_2035_n1610# a_1519_n500# a_545_n2808# a_4615_n500# a_n1319_n1610# a_2293_n2720#
+ a_29_n2808# a_n487_n2808# a_n1577_n2720# a_n2093_n500# a_1519_n1610# a_n4157_n2720#
+ a_1777_n2720#
X0 a_5389_n2720# a_5189_n2808# a_5131_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X1 a_4357_n1610# a_4157_n2808# a_4099_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_n1061_1720# a_n1261_n2808# a_n1319_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_2551_n2720# a_2351_n2808# a_2293_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a_n803_610# a_n1003_n2808# a_n1061_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X5 a_1003_n500# a_803_n2808# a_745_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X6 a_n1835_n2720# a_n2035_n2808# a_n2093_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X7 a_n803_n1610# a_n1003_n2808# a_n1061_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X8 a_745_610# a_545_n2808# a_487_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X9 a_1003_1720# a_803_n2808# a_745_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X10 a_5389_610# a_5189_n2808# a_5131_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X11 a_745_n500# a_545_n2808# a_487_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X12 a_n29_610# a_n229_n2808# a_n287_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X13 a_n3899_610# a_n4099_n2808# a_n4157_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X14 a_1261_n2720# a_1061_n2808# a_1003_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X15 a_745_1720# a_545_n2808# a_487_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X16 a_487_n500# a_287_n2808# a_229_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X17 a_n4931_n2720# a_n5131_n2808# a_n5189_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X18 a_487_1720# a_287_n2808# a_229_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X19 a_n4673_610# a_n4873_n2808# a_n4931_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X20 a_229_n2720# a_29_n2808# a_n29_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X21 a_n545_n2720# a_n745_n2808# a_n803_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X22 a_229_610# a_29_n2808# a_n29_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X23 a_2035_n500# a_1835_n2808# a_1777_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X24 a_4099_n500# a_3899_n2808# a_3841_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X25 a_4099_n2720# a_3899_n2808# a_3841_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X26 a_3067_n1610# a_2867_n2808# a_2809_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X27 a_2035_1720# a_1835_n2808# a_1777_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X28 a_4099_1720# a_3899_n2808# a_3841_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X29 a_n5189_610# a_n5389_n2808# a_n5447_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X30 a_1777_n500# a_1577_n2808# a_1519_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X31 a_4099_610# a_3899_n2808# a_3841_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X32 a_n2609_n500# a_n2809_n2808# a_n2867_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X33 a_3841_n500# a_3641_n2808# a_3583_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X34 a_1777_1720# a_1577_n2808# a_1519_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X35 a_n2609_1720# a_n2809_n2808# a_n2867_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X36 a_3841_1720# a_3641_n2808# a_3583_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X37 a_1519_610# a_1319_n2808# a_1261_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X38 a_3583_n500# a_3383_n2808# a_3325_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X39 a_2809_n1610# a_2609_n2808# a_2551_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X40 a_n4415_n500# a_n4615_n2808# a_n4673_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X41 a_1261_n500# a_1061_n2808# a_1003_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X42 a_1777_n1610# a_1577_n2808# a_1519_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X43 a_n5447_n1610# a_n5647_n2808# a_n5705_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X44 a_3583_1720# a_3383_n2808# a_3325_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X45 a_n3641_n2720# a_n3841_n2808# a_n3899_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X46 a_n4415_1720# a_n4615_n2808# a_n4673_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X47 a_n4157_n500# a_n4357_n2808# a_n4415_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X48 a_1261_1720# a_1061_n2808# a_1003_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X49 a_n3899_n500# a_n4099_n2808# a_n4157_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X50 a_n1835_n500# a_n2035_n2808# a_n2093_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X51 a_n4157_1720# a_n4357_n2808# a_n4415_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X52 a_4873_n1610# a_4673_n2808# a_4615_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X53 a_1519_n1610# a_1319_n2808# a_1261_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X54 a_487_610# a_287_n2808# a_229_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X55 a_n3899_1720# a_n4099_n2808# a_n4157_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X56 a_n1835_1720# a_n2035_n2808# a_n2093_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X57 a_n5189_n2720# a_n5389_n2808# a_n5447_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X58 a_n4157_n1610# a_n4357_n2808# a_n4415_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X59 a_n2351_n2720# a_n2551_n2808# a_n2609_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X60 a_1003_n2720# a_803_n2808# a_745_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X61 a_5647_n2720# a_5447_n2808# a_5389_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X62 a_4615_n1610# a_4415_n2808# a_4357_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X63 a_3583_n1610# a_3383_n2808# a_3325_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X64 a_n545_610# a_n745_n2808# a_n803_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X65 a_2809_610# a_2609_n2808# a_2551_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X66 a_n3899_n2720# a_n4099_n2808# a_n4157_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X67 a_n2867_n1610# a_n3067_n2808# a_n3125_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X68 a_n1319_610# a_n1519_n2808# a_n1577_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X69 a_n1061_n2720# a_n1261_n2808# a_n1319_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X70 a_4357_n2720# a_4157_n2808# a_4099_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X71 a_487_n1610# a_287_n2808# a_229_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X72 a_3325_610# a_3125_n2808# a_3067_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X73 a_3325_n1610# a_3125_n2808# a_3067_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X74 a_2293_n1610# a_2093_n2808# a_2035_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X75 a_n1835_610# a_n2035_n2808# a_n2093_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X76 a_n803_n2720# a_n1003_n2808# a_n1061_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X77 a_1261_610# a_1061_n2808# a_1003_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X78 a_2809_n500# a_2609_n2808# a_2551_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X79 a_n4673_n500# a_n4873_n2808# a_n4931_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X80 a_2809_1720# a_2609_n2808# a_2551_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X81 a_n2609_610# a_n2809_n2808# a_n2867_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X82 a_n287_n1610# a_n487_n2808# a_n545_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X83 a_4615_n500# a_4415_n2808# a_4357_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X84 a_n4673_1720# a_n4873_n2808# a_n4931_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X85 a_4615_610# a_4415_n2808# a_4357_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X86 a_n2351_n500# a_n2551_n2808# a_n2609_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X87 a_4357_n500# a_4157_n2808# a_4099_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X88 a_4615_1720# a_4415_n2808# a_4357_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X89 a_n3125_610# a_n3325_n2808# a_n3383_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X90 a_n2609_n1610# a_n2809_n2808# a_n2867_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X91 a_n2351_1720# a_n2551_n2808# a_n2609_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X92 a_2035_610# a_1835_n2808# a_1777_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X93 a_n2093_n500# a_n2293_n2808# a_n2351_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X94 a_4357_1720# a_4157_n2808# a_4099_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X95 a_229_n500# a_29_n2808# a_n29_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X96 a_n29_n1610# a_n229_n2808# a_n287_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X97 a_n1577_n1610# a_n1777_n2808# a_n1835_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X98 a_n2093_1720# a_n2293_n2808# a_n2351_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X99 a_n29_n500# a_n229_n2808# a_n287_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X100 a_229_1720# a_29_n2808# a_n29_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X101 a_2551_610# a_2351_n2808# a_2293_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X102 a_3067_n2720# a_2867_n2808# a_2809_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X103 a_2035_n1610# a_1835_n2808# a_1777_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X104 a_n29_1720# a_n229_n2808# a_n287_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X105 a_n1061_610# a_n1261_n2808# a_n1319_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X106 a_n1319_n1610# a_n1519_n2808# a_n1577_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X107 a_n4673_n1610# a_n4873_n2808# a_n4931_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X108 a_n287_610# a_n487_n2808# a_n545_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X109 a_2809_n2720# a_2609_n2808# a_2551_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X110 a_5131_n1610# a_4931_n2808# a_4873_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X111 a_1777_n2720# a_1577_n2808# a_1519_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X112 a_n5447_n2720# a_n5647_n2808# a_n5705_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X113 a_n4415_n1610# a_n4615_n2808# a_n4673_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X114 a_n3383_n1610# a_n3583_n2808# a_n3641_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X115 a_n4415_610# a_n4615_n2808# a_n4673_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X116 a_4873_n2720# a_4673_n2808# a_4615_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X117 a_3841_n1610# a_3641_n2808# a_3583_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X118 a_1519_n2720# a_1319_n2808# a_1261_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X119 a_n4931_610# a_n5131_n2808# a_n5189_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X120 a_3841_610# a_3641_n2808# a_3583_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X121 a_n4157_n2720# a_n4357_n2808# a_n4415_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X122 a_n3125_n1610# a_n3325_n2808# a_n3383_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X123 a_n2093_n1610# a_n2293_n2808# a_n2351_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X124 a_n2351_610# a_n2551_n2808# a_n2609_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X125 a_745_n1610# a_545_n2808# a_487_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X126 a_3067_n500# a_2867_n2808# a_2809_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X127 a_4615_n2720# a_4415_n2808# a_4357_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X128 a_5389_n1610# a_5189_n2808# a_5131_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X129 a_3583_n2720# a_3383_n2808# a_3325_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X130 a_2551_n1610# a_2351_n2808# a_2293_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X131 a_5131_n500# a_4931_n2808# a_4873_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X132 a_3067_1720# a_2867_n2808# a_2809_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X133 a_n2867_n2720# a_n3067_n2808# a_n3125_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X134 a_n1835_n1610# a_n2035_n2808# a_n2093_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X135 a_5131_1720# a_4931_n2808# a_4873_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X136 a_4873_n500# a_4673_n2808# a_4615_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X137 a_4357_610# a_4157_n2808# a_4099_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X138 a_3325_n2720# a_3125_n2808# a_3067_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X139 a_487_n2720# a_287_n2808# a_229_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X140 a_4873_1720# a_4673_n2808# a_4615_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X141 a_n1319_n500# a_n1519_n2808# a_n1577_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X142 a_2551_n500# a_2351_n2808# a_2293_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X143 a_n2867_610# a_n3067_n2808# a_n3125_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X144 a_n5447_n500# a_n5647_n2808# a_n5705_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X145 a_2293_n2720# a_2093_n2808# a_2035_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X146 a_1261_n1610# a_1061_n2808# a_1003_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X147 a_n4931_n1610# a_n5131_n2808# a_n5189_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X148 a_1777_610# a_1577_n2808# a_1519_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X149 a_n545_n500# a_n745_n2808# a_n803_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X150 a_2293_n500# a_2093_n2808# a_2035_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X151 a_n1319_1720# a_n1519_n2808# a_n1577_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X152 a_2551_1720# a_2351_n2808# a_2293_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X153 a_n5189_n500# a_n5389_n2808# a_n5447_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X154 a_n5447_1720# a_n5647_n2808# a_n5705_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X155 a_n3125_n500# a_n3325_n2808# a_n3383_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X156 a_n287_n500# a_n487_n2808# a_n545_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X157 a_n545_1720# a_n745_n2808# a_n803_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X158 a_2293_1720# a_2093_n2808# a_2035_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X159 a_2293_610# a_2093_n2808# a_2035_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X160 a_5131_610# a_4931_n2808# a_4873_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X161 a_n2867_n500# a_n3067_n2808# a_n3125_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X162 a_n803_n500# a_n1003_n2808# a_n1061_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X163 a_229_n1610# a_29_n2808# a_n29_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X164 a_n545_n1610# a_n745_n2808# a_n803_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X165 a_n5189_1720# a_n5389_n2808# a_n5447_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X166 a_n3125_1720# a_n3325_n2808# a_n3383_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X167 a_n287_1720# a_n487_n2808# a_n545_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X168 a_n3641_610# a_n3841_n2808# a_n3899_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X169 a_n4931_n500# a_n5131_n2808# a_n5189_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X170 a_n2867_1720# a_n3067_n2808# a_n3125_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X171 a_n803_1720# a_n1003_n2808# a_n1061_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X172 a_n4931_1720# a_n5131_n2808# a_n5189_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X173 a_1003_610# a_803_n2808# a_745_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X174 a_n287_n2720# a_n487_n2808# a_n545_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X175 a_5647_610# a_5447_n2808# a_5389_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X176 a_4099_n1610# a_3899_n2808# a_3841_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X177 a_n4157_610# a_n4357_n2808# a_n4415_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X178 a_3067_610# a_2867_n2808# a_2809_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X179 a_n2609_n2720# a_n2809_n2808# a_n2867_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X180 a_n1577_610# a_n1777_n2808# a_n1835_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X181 a_n29_n2720# a_n229_n2808# a_n287_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X182 a_n1577_n2720# a_n1777_n2808# a_n1835_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X183 a_3583_610# a_3383_n2808# a_3325_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X184 a_2035_n2720# a_1835_n2808# a_1777_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X185 a_n2093_610# a_n2293_n2808# a_n2351_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X186 a_n4673_n2720# a_n4873_n2808# a_n4931_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X187 a_n1319_n2720# a_n1519_n2808# a_n1577_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X188 a_n3641_n1610# a_n3841_n2808# a_n3899_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X189 a_5131_n2720# a_4931_n2808# a_4873_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X190 a_n4415_n2720# a_n4615_n2808# a_n4673_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X191 a_n5189_n1610# a_n5389_n2808# a_n5447_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X192 a_n1577_n500# a_n1777_n2808# a_n1835_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X193 a_n3383_n2720# a_n3583_n2808# a_n3641_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X194 a_n2351_n1610# a_n2551_n2808# a_n2609_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X195 a_n5447_610# a_n5647_n2808# a_n5705_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X196 a_n3641_n500# a_n3841_n2808# a_n3899_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X197 a_1003_n1610# a_803_n2808# a_745_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X198 a_1519_n500# a_1319_n2808# a_1261_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X199 a_5647_n1610# a_5447_n2808# a_5389_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X200 a_5647_n500# a_5447_n2808# a_5389_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X201 a_3841_n2720# a_3641_n2808# a_3583_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X202 a_n1577_1720# a_n1777_n2808# a_n1835_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X203 a_n3383_n500# a_n3583_n2808# a_n3641_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X204 a_n3641_1720# a_n3841_n2808# a_n3899_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X205 a_1519_1720# a_1319_n2808# a_1261_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X206 a_3325_n500# a_3125_n2808# a_3067_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X207 a_n3125_n2720# a_n3325_n2808# a_n3383_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X208 a_5389_n500# a_5189_n2808# a_5131_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X209 a_5647_1720# a_5447_n2808# a_5389_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X210 a_4873_610# a_4673_n2808# a_4615_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X211 a_n3899_n1610# a_n4099_n2808# a_n4157_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X212 a_n3383_1720# a_n3583_n2808# a_n3641_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X213 a_n1061_n500# a_n1261_n2808# a_n1319_n500# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X214 a_n2093_n2720# a_n2293_n2808# a_n2351_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X215 a_n1061_n1610# a_n1261_n2808# a_n1319_n1610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X216 a_3325_1720# a_3125_n2808# a_3067_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X217 a_5389_1720# a_5189_n2808# a_5131_1720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X218 a_n3383_610# a_n3583_n2808# a_n3641_610# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X219 a_745_n2720# a_545_n2808# a_487_n2720# a_n5839_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt Output_OA VDD VOUT VINN VINP VBIAS w_8718_n902# w_7736_n902# VSS w_4240_n902#
XXR1 VSS m1_10706_1822# VOUT sky130_fd_pr__res_high_po_0p69_FJD3D2
Xsky130_fd_pr__nfet_05v0_nvt_FEJX3A_0 VINP VINP w_8718_n902# w_8718_n902# w_8718_n902#
+ m1_9368_n744# w_8718_n902# m1_9368_n744# w_8718_n902# VINP m1_9368_n744# m1_9368_n744#
+ VINP m1_9368_n744# m1_9368_n744# w_8718_n902# VINP w_8718_n902# m1_9368_n744# w_8718_n902#
+ VINP VINP w_8718_n902# w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902# w_8718_n902#
+ VINP VINP w_8718_n902# m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP m1_9368_n744#
+ m1_9368_n744# VINP m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902#
+ VINP VINP w_8718_n902# VINP VINP w_8718_n902# VINP w_8718_n902# w_8718_n902# VINP
+ m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902# m1_9368_n744# w_8718_n902# w_8718_n902#
+ w_8718_n902# VINP w_8718_n902# VINP w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902#
+ w_8718_n902# m1_9368_n744# VINP m1_9368_n744# VINP m1_9368_n744# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
Xsky130_fd_pr__nfet_g5v0d10v5_3WU84W_0 VOUT VSS VSS VOUT VOUT VOUT VSS VSS VOUT VSS
+ w_7736_n902# VOUT VSS VSS VBIAS VOUT VBIAS VSS VOUT VSS VSS VBIAS VOUT VOUT VOUT
+ w_7736_n902# VSS VSS VBIAS VOUT VSS VSS VBIAS VSS VOUT VOUT VSS VSS VSS VSS VSS
+ w_7736_n902# VBIAS VSS VBIAS VBIAS VSS VSS VOUT VSS VSS VBIAS VSS VBIAS VBIAS VBIAS
+ VSS VOUT VOUT VSS VOUT VBIAS VSS VOUT VSS w_7736_n902# VOUT VOUT VSS VSS VOUT VBIAS
+ VSS VSS VSS VOUT VOUT VSS VSS VBIAS VBIAS VSS VSS VSS VOUT VOUT VSS VOUT VOUT VSS
+ VSS VSS VOUT VSS VBIAS w_7736_n902# VOUT VSS VSS VOUT VOUT VOUT VOUT VSS VOUT VBIAS
+ VSS VSS VBIAS VOUT VOUT VBIAS w_7736_n902# VOUT VOUT VOUT VBIAS VOUT VOUT VSS VOUT
+ VBIAS VOUT VBIAS VSS VSS VSS VSS VOUT VSS VBIAS VSS VSS VOUT VOUT VSS VOUT VOUT
+ VSS VSS VOUT VSS VSS VSS VBIAS VOUT VBIAS VOUT VOUT VSS VOUT VSS VSS VOUT VSS VOUT
+ VSS VOUT VBIAS VOUT VOUT VOUT VOUT VBIAS VOUT VSS VSS VBIAS VSS VBIAS VSS VOUT VSS
+ VBIAS VOUT VSS VOUT VSS VSS VSS VSS VOUT w_7736_n902# VSS VSS VSS VSS VSS VSS VBIAS
+ VOUT VBIAS VSS VOUT VOUT VOUT VSS VSS VOUT VOUT VBIAS VSS w_7736_n902# VBIAS VBIAS
+ VOUT VBIAS VOUT VSS VSS VOUT VOUT VSS VSS VOUT VOUT VSS VSS VSS VSS VOUT VSS VOUT
+ w_7736_n902# VSS VSS VOUT VSS VOUT VSS VSS VBIAS VSS VOUT VOUT VBIAS VOUT VOUT VOUT
+ w_7736_n902# VBIAS VOUT VOUT VSS VOUT VSS VOUT VOUT VOUT VOUT VOUT VBIAS VSS VOUT
+ VSS VOUT VSS VSS VSS VBIAS VSS VOUT VOUT VBIAS VBIAS VSS VSS VSS VSS VOUT sky130_fd_pr__nfet_g5v0d10v5_3WU84W
XXM2 VINN w_8718_n902# VINP w_7736_n902# w_7736_n902# w_4240_n902# w_7736_n902# sky130_fd_pr__nfet_01v8_lvt_AJ3MPE
XXM6 m1_9368_n744# m1_4902_n766# m1_9368_n744# VDD m1_4902_n766# m1_4902_n766# VDD
+ m1_4902_n766# m1_4902_n766# m1_4902_n766# VDD sky130_fd_pr__pfet_01v8_lvt_UX3DP3
XXM8 VDD VOUT VDD VOUT VDD VDD VOUT VDD m1_9368_n744# VDD VDD VOUT VOUT m1_9368_n744#
+ VDD VOUT m1_9368_n744# VOUT m1_9368_n744# m1_9368_n744# VOUT VDD m1_9368_n744# m1_9368_n744#
+ VDD VOUT VDD VOUT m1_9368_n744# m1_9368_n744# m1_9368_n744# sky130_fd_pr__pfet_g5v0d10v5_8UL4MK
Xsky130_fd_pr__cap_mim_m3_1_BHK9HY_0 m1_9368_n744# m1_9368_n744# m1_10706_1822# m1_10706_1822#
+ m1_10706_1822# m1_9368_n744# sky130_fd_pr__cap_mim_m3_1_BHK9HY
XXM10 VINN VINN m1_4902_n766# m1_4902_n766# m1_4902_n766# w_4240_n902# m1_4902_n766#
+ w_4240_n902# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902#
+ m1_4902_n766# VINN m1_4902_n766# w_4240_n902# m1_4902_n766# VINN VINN m1_4902_n766#
+ m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# w_4240_n902# VINN VINN m1_4902_n766#
+ w_4240_n902# w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902#
+ w_4240_n902# w_4240_n902# VINN VINN m1_4902_n766# VINN VINN m1_4902_n766# VINN VINN
+ m1_4902_n766# VINN m1_4902_n766# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN
+ VINN m1_4902_n766# w_4240_n902# m1_4902_n766# m1_4902_n766# m1_4902_n766# VINN m1_4902_n766#
+ VINN m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# m1_4902_n766# w_4240_n902#
+ VINN w_4240_n902# VINN w_4240_n902# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_V6AMGK a_n782_n1904# a_9178_n1904# a_13494_1472#
+ a_1376_n1904# a_2704_n1904# a_5194_1472# a_11336_n1904# a_8182_1472# a_6688_n1904#
+ a_n12900_1472# a_546_n1904# a_n10908_n1904# a_n3438_1472# a_10506_1472# a_n6426_1472#
+ a_n2110_1472# a_n12070_n1904# a_n9414_1472# a_n8750_n1904# a_2206_1472# a_12996_1472#
+ a_1708_n1904# a_n10244_1472# a_4696_1472# a_n13232_1472# a_7684_1472# a_48_1472#
+ a_n2442_n1904# a_8182_n1904# a_9510_n1904# a_n11074_n1904# a_n7754_n1904# a_n5928_1472#
+ a_n1612_1472# a_n12402_n1904# a_n4600_1472# a_n8916_1472# a_1708_1472# a_10340_n1904#
+ a_5692_n1904# a_n9248_n1904# a_3202_n1904# a_n12734_1472# a_n1446_n1904# a_n13896_n1904#
+ a_2870_1472# a_7186_n1904# a_8514_n1904# a_n10078_n1904# a_n6758_n1904# a_712_1472#
+ a_13328_1472# a_n11406_n1904# a_12000_1472# a_n9248_1472# a_n284_n1904# a_4696_n1904#
+ a_n948_1472# a_5028_1472# a_8016_1472# a_n10078_1472# a_2206_n1904# a_n13066_1472#
+ a_6190_1472# a_7518_n1904# a_n1446_1472# a_n4434_1472# a_11502_1472# a_n8252_n1904#
+ a_n616_n1904# a_n7422_1472# a_3202_1472# a_7518_1472# a_13992_1472# a_6190_n1904#
+ a_n12568_1472# a_n5762_n1904# a_n10410_n1904# a_n11240_1472# a_5692_1472# a_8680_1472#
+ a_546_1472# a_9012_n1904# a_n7256_n1904# a_13660_n1904# a_n3936_1472# a_1210_n1904#
+ a_n6924_1472# a_5194_n1904# a_n9912_1472# a_2704_1472# a_6522_n1904# a_n4766_n1904#
+ a_n10742_1472# a_n13398_n1904# a_n13730_1472# a_8016_n1904# a_12664_n1904# a_n4268_1472#
+ a_11336_1472# a_n7256_1472# a_4198_n1904# a_5526_n1904# a_3036_1472# a_14158_n1904#
+ a_6024_1472# a_9012_1472# a_n11074_1472# a_n6260_n1904# a_n14062_1472# a_11668_n1904#
+ a_878_n1904# a_10838_1472# a_n3770_n1904# a_n118_n1904# a_n6758_1472# a_n2442_1472#
+ a_13826_1472# a_n9746_1472# a_n5430_1472# a_2538_1472# a_n13730_n1904# a_1210_1472#
+ a_5526_1472# a_7020_n1904# a_n5264_n1904# a_8514_1472# a_n10576_1472# a_n13564_1472#
+ a_4530_n1904# a_n2774_n1904# a_14158_1472# a_13162_n1904# a_n1944_1472# a_9842_n1904#
+ a_n4932_1472# a_n12734_n1904# a_6024_n1904# a_n7920_1472# a_n4268_n1904# a_n450_1472#
+ a_10672_n1904# a_3700_1472# a_n14228_n1904# a_3534_n1904# a_n1778_n1904# a_12166_n1904#
+ a_n2276_1472# a_8846_n1904# a_12332_1472# a_n5264_1472# a_n11738_n1904# a_5028_n1904#
+ a_n8252_1472# a_1044_1472# a_4032_1472# a_8348_1472# a_n9580_n1904# a_7020_1472#
+ a_n13398_1472# a_2538_n1904# a_n12070_1472# a_n14358_n2034# a_n3272_n1904# a_n1778_1472#
+ a_n4766_1472# a_n4600_n1904# a_11834_1472# a_n7754_1472# a_n8584_n1904# a_n948_n1904#
+ a_n284_1472# a_n13232_n1904# a_n9912_n1904# a_3534_1472# a_11170_n1904# a_6522_1472#
+ a_380_n1904# a_7850_n1904# a_9510_1472# a_n11572_1472# a_n10742_n1904# a_4032_n1904#
+ a_n2276_n1904# a_878_1472# a_n5098_1472# a_n3604_n1904# a_12166_1472# a_9344_n1904#
+ a_n7588_n1904# a_n8086_1472# a_13992_n1904# a_n12236_n1904# a_n8916_n1904# a_n2940_1472#
+ a_1542_n1904# a_10174_n1904# a_11502_n1904# a_6854_n1904# a_712_n1904# a_3036_n1904#
+ a_n2608_n1904# a_8348_n1904# a_12996_n1904# a_11668_1472# a_n3272_1472# a_10340_1472#
+ a_n7588_1472# a_n6260_1472# a_3368_1472# a_10506_n1904# a_n9082_n1904# a_5858_n1904#
+ a_2040_1472# a_6356_1472# a_9344_1472# a_n1280_n1904# a_n6592_n1904# a_n11240_n1904#
+ a_n7920_n1904# a_n118_1472# a_n4102_n1904# a_n2774_1472# a_n8086_n1904# a_n5762_1472#
+ a_12830_1472# a_n9414_n1904# a_2040_n1904# a_n8750_1472# a_n11406_1472# a_1542_1472#
+ a_5858_1472# a_n1612_n1904# a_12000_n1904# a_4530_1472# a_8846_1472# a_7352_n1904#
+ a_n5596_n1904# a_n13896_1472# a_n10244_n1904# a_n6924_n1904# a_n3106_n1904# a_n450_n1904#
+ a_10174_1472# a_4862_n1904# a_13494_n1904# a_n6094_1472# a_13162_1472# a_n8418_n1904#
+ a_1044_n1904# a_n9082_1472# a_11004_n1904# a_n10908_1472# a_9178_1472# a_n782_1472#
+ a_6356_n1904# a_214_n1904# a_n5928_n1904# a_n3106_1472# a_n7090_n1904# a_3866_n1904#
+ a_12498_n1904# a_13826_n1904# a_n5596_1472# a_n1280_1472# a_12664_1472# a_10008_n1904#
+ a_n8584_1472# a_1376_1472# a_n14228_1472# a_4364_1472# a_7352_1472# a_n2110_n1904#
+ a_n6094_n1904# a_n7422_n1904# a_n2608_1472# a_380_1472# a_5360_n1904# a_n4932_n1904#
+ a_n3770_1472# a_n1114_n1904# a_n13564_n1904# a_3866_1472# a_n12402_1472# a_n5098_n1904#
+ a_2870_n1904# a_6854_1472# a_n6426_n1904# a_9842_1472# a_12830_n1904# a_10008_1472#
+ a_4364_n1904# a_12498_1472# a_n3936_n1904# a_n616_1472# a_11170_1472# a_9676_n1904#
+ a_n7090_1472# a_n12568_n1904# a_4198_1472# a_1874_n1904# a_7186_1472# a_n11904_1472#
+ a_11834_n1904# a_n1114_1472# a_3368_n1904# a_n4102_1472# a_n8418_1472# a_13328_n1904#
+ a_48_n1904# a_10672_1472# a_n6592_1472# a_13660_1472# a_n5430_n1904# a_n9580_1472#
+ a_n12236_1472# a_6688_1472# a_10838_n1904# a_2372_1472# a_n14062_n1904# a_5360_1472#
+ a_9676_1472# a_214_1472# a_n2940_n1904# a_8680_n1904# a_n3604_1472# a_n11572_n1904#
+ a_n12900_n1904# a_n4434_n1904# a_n11738_1472# a_n13066_n1904# a_n9746_n1904# a_1874_1472#
+ a_2372_n1904# a_n10410_1472# a_4862_1472# a_3700_n1904# a_n1944_n1904# a_12332_n1904#
+ a_7850_1472# a_7684_n1904# a_n10576_n1904# a_11004_1472# a_n11904_n1904# a_n3438_n1904#
X0 a_8016_1472# a_8016_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X1 a_n616_1472# a_n616_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X2 a_3368_1472# a_3368_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X3 a_1044_1472# a_1044_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X4 a_n6924_1472# a_n6924_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X5 a_n9746_1472# a_n9746_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X6 a_n7422_1472# a_n7422_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X7 a_546_1472# a_546_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X8 a_380_1472# a_380_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X9 a_n13896_1472# a_n13896_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X10 a_n11738_1472# a_n11738_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X11 a_n11572_1472# a_n11572_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X12 a_n2940_1472# a_n2940_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X13 a_n2774_1472# a_n2774_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X14 a_n12236_1472# a_n12236_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X15 a_13826_1472# a_13826_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X16 a_11502_1472# a_11502_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X17 a_n3438_1472# a_n3438_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X18 a_13660_1472# a_13660_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X19 a_7850_1472# a_7850_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X20 a_n1114_1472# a_n1114_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X21 a_n5596_1472# a_n5596_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X22 a_n3272_1472# a_n3272_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X23 a_12000_1472# a_12000_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X24 a_8514_1472# a_8514_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X25 a_n6260_1472# a_n6260_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X26 a_n6094_1472# a_n6094_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X27 a_3866_1472# a_3866_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X28 a_1708_1472# a_1708_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X29 a_1542_1472# a_1542_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X30 a_9012_1472# a_9012_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X31 a_12498_1472# a_12498_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X32 a_10174_1472# a_10174_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X33 a_6688_1472# a_6688_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X34 a_4364_1472# a_4364_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X35 a_2206_1472# a_2206_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X36 a_2040_1472# a_2040_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X37 a_5028_1472# a_5028_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X38 a_7186_1472# a_7186_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X39 a_n12734_1472# a_n12734_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X40 a_n450_1472# a_n450_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X41 a_n3936_1472# a_n3936_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X42 a_n284_1472# a_n284_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X43 a_n1612_1472# a_n1612_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X44 a_n13232_1472# a_n13232_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X45 a_n6758_1472# a_n6758_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X46 a_n4434_1472# a_n4434_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X47 a_48_1472# a_48_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X48 a_n6592_1472# a_n6592_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X49 a_9510_1472# a_9510_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X50 a_n9580_1472# a_n9580_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X51 a_n7256_1472# a_n7256_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X52 a_10838_1472# a_10838_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X53 a_2704_1472# a_2704_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X54 a_12996_1472# a_12996_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X55 a_10672_1472# a_10672_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X56 a_4862_1472# a_4862_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X57 a_n12070_1472# a_n12070_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X58 a_13494_1472# a_13494_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X59 a_11336_1472# a_11336_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X60 a_7684_1472# a_7684_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X61 a_5526_1472# a_5526_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X62 a_5360_1472# a_5360_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X63 a_3202_1472# a_3202_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X64 a_11170_1472# a_11170_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X65 a_14158_1472# a_14158_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X66 a_8348_1472# a_8348_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X67 a_8182_1472# a_8182_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X68 a_6024_1472# a_6024_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X69 a_n782_1472# a_n782_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X70 a_n948_1472# a_n948_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X71 a_1376_1472# a_1376_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X72 a_n4932_1472# a_n4932_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X73 a_4198_1472# a_4198_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X74 a_n7920_1472# a_n7920_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X75 a_n7754_1472# a_n7754_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X76 a_878_1472# a_878_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X77 a_n8418_1472# a_n8418_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X78 a_n8252_1472# a_n8252_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X79 a_n10410_1472# a_n10410_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X80 a_n12568_1472# a_n12568_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X81 a_n10244_1472# a_n10244_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X82 a_11834_1472# a_11834_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X83 a_3700_1472# a_3700_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X84 a_n3770_1472# a_n3770_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X85 a_13992_1472# a_13992_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X86 a_n1446_1472# a_n1446_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X87 a_n13066_1472# a_n13066_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X88 a_n2110_1472# a_n2110_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X89 a_12332_1472# a_12332_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X90 a_8846_1472# a_8846_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X91 a_6522_1472# a_6522_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X92 a_n4268_1472# a_n4268_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X93 a_8680_1472# a_8680_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X94 a_1874_1472# a_1874_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X95 a_9344_1472# a_9344_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X96 a_7020_1472# a_7020_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X97 a_n7090_1472# a_n7090_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X98 a_4696_1472# a_4696_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X99 a_2538_1472# a_2538_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X100 a_2372_1472# a_2372_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X101 a_5194_1472# a_5194_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X102 a_3036_1472# a_3036_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X103 a_n8916_1472# a_n8916_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X104 a_n10908_1472# a_n10908_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X105 a_n10742_1472# a_n10742_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X106 a_n9414_1472# a_n9414_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X107 a_n1944_1472# a_n1944_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X108 a_n13730_1472# a_n13730_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X109 a_n11406_1472# a_n11406_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X110 a_214_1472# a_214_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X111 a_n13564_1472# a_n13564_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X112 a_n4766_1472# a_n4766_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X113 a_n2608_1472# a_n2608_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X114 a_12830_1472# a_12830_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X115 a_n2442_1472# a_n2442_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X116 a_n14228_1472# a_n14228_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X117 a_n14062_1472# a_n14062_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X118 a_9842_1472# a_9842_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X119 a_n7588_1472# a_n7588_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X120 a_n5430_1472# a_n5430_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X121 a_n5264_1472# a_n5264_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X122 a_n3106_1472# a_n3106_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X123 a_2870_1472# a_2870_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X124 a_n8086_1472# a_n8086_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X125 a_n10078_1472# a_n10078_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X126 a_11668_1472# a_11668_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X127 a_5858_1472# a_5858_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X128 a_3534_1472# a_3534_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X129 a_1210_1472# a_1210_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X130 a_5692_1472# a_5692_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X131 a_n1280_1472# a_n1280_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X132 a_10008_1472# a_10008_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X133 a_12166_1472# a_12166_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X134 a_6356_1472# a_6356_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X135 a_4032_1472# a_4032_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X136 a_6190_1472# a_6190_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X137 a_n9912_1472# a_n9912_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X138 a_712_1472# a_712_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X139 a_n11904_1472# a_n11904_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X140 a_9178_1472# a_9178_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X141 a_n12402_1472# a_n12402_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X142 a_n118_1472# a_n118_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X143 a_n5928_1472# a_n5928_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X144 a_n3604_1472# a_n3604_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X145 a_n5762_1472# a_n5762_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X146 a_n8750_1472# a_n8750_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X147 a_n6426_1472# a_n6426_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X148 a_n4102_1472# a_n4102_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X149 a_n8584_1472# a_n8584_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X150 a_n12900_1472# a_n12900_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X151 a_n10576_1472# a_n10576_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X152 a_n1778_1472# a_n1778_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X153 a_n9248_1472# a_n9248_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X154 a_n11240_1472# a_n11240_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X155 a_n9082_1472# a_n9082_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X156 a_n13398_1472# a_n13398_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X157 a_n11074_1472# a_n11074_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X158 a_12664_1472# a_12664_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X159 a_10506_1472# a_10506_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X160 a_10340_1472# a_10340_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X161 a_6854_1472# a_6854_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X162 a_4530_1472# a_4530_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X163 a_n4600_1472# a_n4600_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X164 a_n2276_1472# a_n2276_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X165 a_13328_1472# a_13328_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X166 a_13162_1472# a_13162_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X167 a_11004_1472# a_11004_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X168 a_9676_1472# a_9676_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X169 a_7518_1472# a_7518_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X170 a_7352_1472# a_7352_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
X171 a_n5098_1472# a_n5098_n1904# a_n14358_n2034# sky130_fd_pr__res_xhigh_po_0p35 l=14.88
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_S4N9LQ a_1708_1984# a_n1778_n2416# a_712_1984#
+ a_n948_1984# a_2538_n2416# a_n1446_1984# a_n948_n2416# a_380_n2416# a_546_1984#
+ a_n2276_n2416# a_1542_n2416# a_712_n2416# a_n2608_n2416# a_n1280_n2416# a_n2442_1984#
+ a_2538_1984# a_1210_1984# a_2040_n2416# a_n1612_n2416# a_n1944_1984# a_n450_n2416#
+ a_1044_n2416# a_n450_1984# a_214_n2416# a_n2276_1984# a_1044_1984# a_n2110_n2416#
+ a_n1778_1984# a_n284_1984# a_n1114_n2416# a_878_1984# a_1874_n2416# a_48_n2416#
+ a_2040_1984# a_n118_1984# a_n2738_n2546# a_1542_1984# a_2372_n2416# a_n1944_n2416#
+ a_n782_n2416# a_n782_1984# a_1376_n2416# a_546_n2416# a_n1280_1984# a_1376_1984#
+ a_1708_n2416# a_n2442_n2416# a_n2608_1984# a_380_1984# a_n1446_n2416# a_n616_1984#
+ a_n284_n2416# a_2206_n2416# a_n1114_1984# a_n616_n2416# a_2372_1984# a_214_1984#
+ a_1210_n2416# a_1874_1984# a_878_n2416# a_n2110_1984# a_n118_n2416# a_2206_1984#
+ a_48_1984# a_n1612_1984#
X0 a_2040_1984# a_2040_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X1 a_2206_1984# a_2206_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X2 a_n450_1984# a_n450_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X3 a_n284_1984# a_n284_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X4 a_n1612_1984# a_n1612_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X5 a_48_1984# a_48_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X6 a_n948_1984# a_n948_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X7 a_n782_1984# a_n782_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X8 a_1376_1984# a_1376_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X9 a_878_1984# a_878_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X10 a_n1446_1984# a_n1446_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X11 a_n2110_1984# a_n2110_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X12 a_1874_1984# a_1874_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X13 a_2372_1984# a_2372_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X14 a_2538_1984# a_2538_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X15 a_n1944_1984# a_n1944_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X16 a_n2608_1984# a_n2608_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X17 a_n2442_1984# a_n2442_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X18 a_214_1984# a_214_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X19 a_n1280_1984# a_n1280_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X20 a_1210_1984# a_1210_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X21 a_712_1984# a_712_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X22 a_n118_1984# a_n118_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X23 a_n2276_1984# a_n2276_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X24 a_n1778_1984# a_n1778_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X25 a_n616_1984# a_n616_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X26 a_1044_1984# a_1044_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X27 a_546_1984# a_546_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X28 a_380_1984# a_380_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X29 a_n1114_1984# a_n1114_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X30 a_1542_1984# a_1542_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X31 a_1708_1984# a_1708_n2416# a_n2738_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
.ends

.subckt Parallel_10B_Block2 V6 V5 V8 V9 V7 VO1 VOUT V4 V3 V2 V1 V0 VCM w_8036_n6718#
+ VBIAS w_8040_12750# w_3572_3030# w_3570_n6718# w_8038_3030# w_3574_12750# DVDD w_7054_n6718#
+ w_7056_3030# DVSS AVSS AVDD w_7058_12750#
Xx1 V8 DVDD x7/VINN VCM x1/R2RIN x13/R2RIN AVSS DVSS AVDD Universal_R_2R_Block2
Xx2 V5 DVDD x7/VINN VCM x6/VOUT x5/R2RIN AVSS DVSS AVDD Universal_R_2R_Block2
Xx3 V2 DVDD x7/VINN VCM x3/R2RIN x3/R2ROUT AVSS DVSS AVDD Universal_R_2R_Block2
Xx4 V0 DVDD x7/VINN VCM x8/VOUT x4/R2ROUT AVSS DVSS AVDD Universal_R_2R_Block2
Xx5 V6 DVDD x7/VINN VCM x5/R2RIN x5/R2ROUT AVSS DVSS AVDD Universal_R_2R_Block2
Xx6 AVDD x6/VOUT x6/VINN VCM VBIAS w_3574_12750# w_7058_12750# AVSS w_8040_12750#
+ x1_x32_OA
Xx7 AVDD VOUT x7/VINN VCM VBIAS w_3570_n6718# w_7054_n6718# AVSS w_8036_n6718# Output_OA
Xx8 AVDD x8/VOUT x8/VINN VCM VBIAS w_3572_3030# w_7056_3030# AVSS w_8038_3030# x1_x32_OA
Xx9 V4 DVDD x7/VINN VCM x9/R2RIN x9/R2ROUT AVSS DVSS AVDD Universal_R_2R_Block2
Xsky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_0 m1_13604_18506# VCM m1_13272_18506# m1_12290_20904#
+ AVSS m1_12940_18506# m1_13272_18506# m1_13438_20902# x13/R2ROUT m1_13604_18506#
+ m1_13438_20902# x6/VOUT m1_12940_18506# sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP
Xsky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_1 m1_10646_18508# m1_10146_20906# m1_10314_18508#
+ x9/R2ROUT AVSS m1_9982_18508# m1_10314_18508# VCM VO1 m1_10646_18508# x8/VINN m1_10146_20906#
+ m1_9982_18508# sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP
Xsky130_fd_pr__res_xhigh_po_0p35_Q2LWZP_2 m1_12122_18506# m1_11626_20906# m1_11790_18506#
+ VO1 AVSS m1_11458_18506# m1_11790_18506# x6/VINN m1_12290_20904# m1_12122_18506#
+ x6/VINN m1_11626_20906# m1_11458_18506# sky130_fd_pr__res_xhigh_po_0p35_Q2LWZP
Xx10 V3 DVDD x7/VINN VCM x3/R2ROUT x9/R2RIN AVSS DVSS AVDD Universal_R_2R_Block2
Xx11 V1 DVDD x7/VINN VCM x4/R2ROUT x3/R2RIN AVSS DVSS AVDD Universal_R_2R_Block2
Xx12 V7 DVDD x7/VINN VCM x5/R2ROUT x1/R2RIN AVSS DVSS AVDD Universal_R_2R_Block2
Xx13 V9 DVDD x7/VINN VCM x13/R2RIN x13/R2ROUT AVSS DVSS AVDD Universal_R_2R_Block2
Xsky130_fd_pr__res_xhigh_po_0p35_V6AMGK_0 m1_13942_n11110# m1_23902_n11110# m1_28384_n7734#
+ m1_16266_n11110# m1_17594_n11110# m1_20084_n7734# m1_26226_n11110# m1_23072_n7734#
+ m1_21578_n11110# m1_1824_n7734# m1_15270_n11110# m1_3982_n11110# m1_11452_n7734#
+ m1_25396_n7734# m1_8464_n7734# m1_12780_n7734# m1_2654_n11110# m1_5476_n7734# m1_5974_n11110#
+ m1_17096_n7734# m1_27720_n7734# m1_16598_n11110# m1_4480_n7734# m1_19420_n7734#
+ m1_1492_n7734# m1_22408_n7734# x7/VINN m1_12282_n11110# m1_22906_n11110# m1_24234_n11110#
+ m1_3650_n11110# m1_6970_n11110# m1_8796_n7734# m1_13112_n7734# m1_2322_n11110# m1_10124_n7734#
+ m1_5808_n7734# m1_16432_n7734# m1_25230_n11110# m1_20582_n11110# m1_5642_n11110#
+ m1_17926_n11110# m1_2156_n7734# m1_13278_n11110# m1_994_n11110# m1_17760_n7734#
+ m1_21910_n11110# m1_23238_n11110# m1_4646_n11110# m1_7966_n11110# m1_15436_n7734#
+ m1_28052_n7734# m1_3318_n11110# m1_26724_n7734# m1_5476_n7734# m1_14606_n11110#
+ m1_19586_n11110# m1_13776_n7734# m1_19752_n7734# m1_22740_n7734# m1_4812_n7734#
+ m1_16930_n11110# m1_1824_n7734# m1_21080_n7734# m1_22242_n11110# m1_13444_n7734#
+ m1_10456_n7734# m1_26392_n7734# m1_6638_n11110# m1_14274_n11110# m1_7468_n7734#
+ m1_18092_n7734# m1_22408_n7734# m1_28716_n7734# m1_20914_n11110# m1_2156_n7734#
+ m1_8962_n11110# m1_4314_n11110# m1_3484_n7734# m1_20416_n7734# m1_23404_n7734# m1_15436_n7734#
+ m1_23902_n11110# m1_7634_n11110# m1_28550_n11110# m1_10788_n7734# m1_15934_n11110#
+ m1_7800_n7734# m1_19918_n11110# m1_4812_n7734# m1_17428_n7734# m1_21246_n11110#
+ m1_9958_n11110# m1_4148_n7734# m1_1326_n11110# m1_1160_n7734# m1_22906_n11110# m1_27554_n11110#
+ m1_10456_n7734# m1_26060_n7734# m1_7468_n7734# m1_18922_n11110# m1_20250_n11110#
+ m1_17760_n7734# m1_28882_n11110# m1_20748_n7734# m1_23736_n7734# m1_3816_n7734#
+ m1_8630_n11110# m1_828_n7734# m1_26558_n11110# m1_15602_n11110# m1_25728_n7734#
+ m1_10954_n11110# m1_14606_n11110# m1_8132_n7734# m1_12448_n7734# m1_28716_n7734#
+ m1_5144_n7734# m1_9460_n7734# m1_17428_n7734# m1_994_n11110# m1_16100_n7734# m1_20416_n7734#
+ m1_21910_n11110# m1_9626_n11110# m1_23404_n7734# m1_4148_n7734# m1_1160_n7734# m1_19254_n11110#
+ m1_11950_n11110# VOUT m1_27886_n11110# m1_12780_n7734# m1_24566_n11110# m1_9792_n7734#
+ m1_1990_n11110# m1_20914_n11110# m1_6804_n7734# m1_10622_n11110# m1_14440_n7734#
+ m1_25562_n11110# m1_18424_n7734# m1_662_n11110# m1_18258_n11110# m1_12946_n11110#
+ m1_26890_n11110# m1_12448_n7734# m1_23570_n11110# m1_27056_n7734# m1_9460_n7734#
+ m1_2986_n11110# m1_19918_n11110# m1_6472_n7734# m1_15768_n7734# m1_18756_n7734#
+ m1_23072_n7734# m1_5310_n11110# m1_21744_n7734# m1_1492_n7734# m1_17262_n11110#
+ m1_2820_n7734# AVSS m1_11618_n11110# m1_13112_n7734# m1_10124_n7734# m1_10290_n11110#
+ m1_26724_n7734# m1_7136_n7734# m1_6306_n11110# m1_13942_n11110# m1_14440_n7734#
+ m1_1658_n11110# m1_4978_n11110# m1_18424_n7734# m1_25894_n11110# m1_21412_n7734#
+ m1_15270_n11110# m1_22574_n11110# m1_24400_n7734# m1_3152_n7734# m1_3982_n11110#
+ m1_18922_n11110# m1_12614_n11110# m1_15768_n7734# m1_9792_n7734# m1_11286_n11110#
+ m1_27056_n7734# m1_24234_n11110# m1_7302_n11110# m1_6804_n7734# m1_28882_n11110#
+ m1_2654_n11110# m1_5974_n11110# m1_11784_n7734# m1_16266_n11110# m1_24898_n11110#
+ m1_26226_n11110# m1_21578_n11110# m1_15602_n11110# m1_17926_n11110# m1_12282_n11110#
+ m1_23238_n11110# m1_27886_n11110# m1_26392_n7734# m1_11452_n7734# m1_25064_n7734#
+ m1_7136_n7734# m1_8464_n7734# m1_18092_n7734# m1_25230_n11110# m1_5642_n11110# m1_20582_n11110#
+ m1_16764_n7734# m1_21080_n7734# m1_24068_n7734# m1_13610_n11110# m1_8298_n11110#
+ m1_3650_n11110# m1_6970_n11110# x7/VINN m1_10622_n11110# m1_12116_n7734# m1_6638_n11110#
+ m1_9128_n7734# m1_27720_n7734# m1_5310_n11110# m1_16930_n11110# m1_6140_n7734# m1_3484_n7734#
+ m1_16432_n7734# m1_20748_n7734# m1_13278_n11110# m1_26890_n11110# m1_19420_n7734#
+ m1_23736_n7734# m1_22242_n11110# m1_9294_n11110# m1_828_n7734# m1_4646_n11110# m1_7966_n11110#
+ m1_11618_n11110# m1_14274_n11110# m1_25064_n7734# m1_19586_n11110# m1_28218_n11110#
+ m1_8796_n7734# m1_28052_n7734# m1_6306_n11110# m1_15934_n11110# m1_5808_n7734# m1_25894_n11110#
+ m1_3816_n7734# m1_24068_n7734# m1_14108_n7734# m1_21246_n11110# m1_14938_n11110#
+ m1_8962_n11110# m1_11784_n7734# m1_7634_n11110# m1_18590_n11110# m1_27222_n11110#
+ m1_28550_n11110# m1_9128_n7734# m1_13444_n7734# m1_27388_n7734# m1_24898_n11110#
+ m1_6140_n7734# m1_16100_n7734# x6/VOUT m1_19088_n7734# m1_22076_n7734# m1_12614_n11110#
+ m1_8630_n11110# m1_7302_n11110# m1_12116_n7734# m1_15104_n7734# m1_20250_n11110#
+ m1_9958_n11110# m1_11120_n7734# m1_13610_n11110# m1_1326_n11110# m1_18756_n7734#
+ m1_2488_n7734# m1_9626_n11110# m1_17594_n11110# m1_21744_n7734# m1_8298_n11110#
+ m1_24732_n7734# m1_27554_n11110# m1_24732_n7734# m1_19254_n11110# m1_27388_n7734#
+ m1_10954_n11110# m1_14108_n7734# m1_26060_n7734# m1_24566_n11110# m1_7800_n7734#
+ m1_2322_n11110# m1_19088_n7734# m1_16598_n11110# m1_22076_n7734# m1_2820_n7734#
+ m1_26558_n11110# m1_13776_n7734# m1_18258_n11110# m1_10788_n7734# m1_6472_n7734#
+ m1_28218_n11110# m1_14938_n11110# m1_25396_n7734# m1_8132_n7734# m1_28384_n7734#
+ m1_9294_n11110# m1_5144_n7734# m1_2488_n7734# m1_21412_n7734# m1_25562_n11110# m1_17096_n7734#
+ m1_662_n11110# m1_20084_n7734# m1_24400_n7734# m1_15104_n7734# m1_11950_n11110#
+ m1_23570_n11110# m1_11120_n7734# m1_3318_n11110# m1_1990_n11110# m1_10290_n11110#
+ m1_3152_n7734# m1_1658_n11110# m1_4978_n11110# m1_16764_n7734# m1_17262_n11110#
+ m1_4480_n7734# m1_19752_n7734# m1_18590_n11110# m1_12946_n11110# m1_27222_n11110#
+ m1_22740_n7734# m1_22574_n11110# m1_4314_n11110# m1_25728_n7734# m1_2986_n11110#
+ m1_11286_n11110# sky130_fd_pr__res_xhigh_po_0p35_V6AMGK
Xsky130_fd_pr__res_xhigh_po_0p35_S4N9LQ_0 m1_14152_11224# m1_10666_6824# m1_13156_11224#
+ m1_11496_11224# x8/VINN m1_10832_11224# m1_11330_6824# m1_12658_6824# m1_12824_11224#
+ m1_10002_6824# m1_13986_6824# m1_12990_6824# x8/VOUT m1_10998_6824# m1_9836_11224#
+ m1_14816_11224# m1_13488_11224# m1_14318_6824# m1_10666_6824# m1_10500_11224# m1_11994_6824#
+ m1_13322_6824# m1_11828_11224# m1_12658_6824# m1_10168_11224# m1_13488_11224# m1_10334_6824#
+ m1_10500_11224# m1_12160_11224# m1_11330_6824# m1_13156_11224# m1_14318_6824# m1_12326_6824#
+ m1_14484_11224# m1_12160_11224# AVSS m1_13820_11224# m1_14650_6824# m1_10334_6824#
+ m1_11662_6824# m1_11496_11224# m1_13654_6824# m1_12990_6824# m1_11164_11224# m1_13820_11224#
+ m1_13986_6824# m1_10002_6824# m1_9836_11224# m1_12824_11224# m1_10998_6824# m1_11828_11224#
+ m1_11994_6824# m1_14650_6824# m1_11164_11224# m1_11662_6824# m1_14816_11224# m1_12492_11224#
+ m1_13654_6824# m1_14152_11224# m1_13322_6824# m1_10168_11224# m1_12326_6824# m1_14484_11224#
+ m1_12492_11224# m1_10832_11224# sky130_fd_pr__res_xhigh_po_0p35_S4N9LQ
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_7WHXCK a_n29_n2720# a_487_n1610# a_n287_610#
+ a_229_n2720# a_n803_n2720# a_n287_n1610# a_n287_n500# a_229_1720# a_n745_n2808#
+ a_745_n500# a_n545_1720# a_745_n1610# a_n545_n1610# a_n803_610# a_229_n500# a_n29_n1610#
+ a_n29_1720# a_n229_n2808# a_n803_n1610# a_487_1720# a_487_n2720# a_229_n1610# a_n545_n500#
+ a_745_610# a_n287_n2720# a_229_610# a_n803_1720# a_n545_610# a_287_n2808# a_745_n2720#
+ a_n545_n2720# a_n29_n500# a_487_n500# a_n287_1720# a_487_610# a_n937_n2942# a_n29_610#
+ a_745_1720# a_n803_n500# a_545_n2808# a_29_n2808# a_n487_n2808#
X0 a_n29_610# a_n229_n2808# a_n287_610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X1 a_745_610# a_545_n2808# a_487_610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X2 a_745_n500# a_545_n2808# a_487_n500# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X3 a_487_1720# a_287_n2808# a_229_1720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a_745_1720# a_545_n2808# a_487_1720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X5 a_487_n500# a_287_n2808# a_229_n500# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X6 a_229_610# a_29_n2808# a_n29_610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X7 a_n545_n2720# a_n745_n2808# a_n803_n2720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X8 a_229_n2720# a_29_n2808# a_n29_n2720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X9 a_487_610# a_287_n2808# a_229_610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X10 a_n545_610# a_n745_n2808# a_n803_610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X11 a_487_n1610# a_287_n2808# a_229_n1610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X12 a_n287_n1610# a_n487_n2808# a_n545_n1610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X13 a_229_n500# a_29_n2808# a_n29_n500# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X14 a_n29_n1610# a_n229_n2808# a_n287_n1610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X15 a_229_1720# a_29_n2808# a_n29_1720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X16 a_n29_n500# a_n229_n2808# a_n287_n500# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X17 a_n29_1720# a_n229_n2808# a_n287_1720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X18 a_n287_610# a_n487_n2808# a_n545_610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X19 a_745_n1610# a_545_n2808# a_487_n1610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X20 a_487_n2720# a_287_n2808# a_229_n2720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X21 a_n545_1720# a_n745_n2808# a_n803_1720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X22 a_n545_n500# a_n745_n2808# a_n803_n500# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X23 a_n287_n500# a_n487_n2808# a_n545_n500# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X24 a_n287_1720# a_n487_n2808# a_n545_1720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X25 a_n545_n1610# a_n745_n2808# a_n803_n1610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X26 a_229_n1610# a_29_n2808# a_n29_n1610# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X27 a_n287_n2720# a_n487_n2808# a_n545_n2720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X28 a_n29_n2720# a_n229_n2808# a_n287_n2720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X29 a_745_n2720# a_545_n2808# a_487_n2720# a_n937_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt Input_Stage_OA1 VDD VOUT VINN VINP VBIAS w_8718_n902# w_7736_n902# VSS w_4240_n902#
XXR1 VSS m1_10706_1822# VOUT sky130_fd_pr__res_high_po_0p69_FJD3D2
Xsky130_fd_pr__nfet_05v0_nvt_FEJX3A_0 VINP VINP w_8718_n902# w_8718_n902# w_8718_n902#
+ m1_9368_n744# w_8718_n902# m1_9368_n744# w_8718_n902# VINP m1_9368_n744# m1_9368_n744#
+ VINP m1_9368_n744# m1_9368_n744# w_8718_n902# VINP w_8718_n902# m1_9368_n744# w_8718_n902#
+ VINP VINP w_8718_n902# w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902# w_8718_n902#
+ VINP VINP w_8718_n902# m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP m1_9368_n744#
+ m1_9368_n744# VINP m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902#
+ VINP VINP w_8718_n902# VINP VINP w_8718_n902# VINP w_8718_n902# w_8718_n902# VINP
+ m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902# m1_9368_n744# w_8718_n902# w_8718_n902#
+ w_8718_n902# VINP w_8718_n902# VINP w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902#
+ w_8718_n902# m1_9368_n744# VINP m1_9368_n744# VINP m1_9368_n744# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
XXM2 VINN w_8718_n902# VINP w_7736_n902# w_7736_n902# w_4240_n902# w_7736_n902# sky130_fd_pr__nfet_01v8_lvt_AJ3MPE
XXM6 m1_9368_n744# m1_4902_n766# m1_9368_n744# VDD m1_4902_n766# m1_4902_n766# VDD
+ m1_4902_n766# m1_4902_n766# m1_4902_n766# VDD sky130_fd_pr__pfet_01v8_lvt_UX3DP3
XXM8 VDD VOUT VDD VOUT VDD VDD VOUT VDD m1_9368_n744# VDD VDD VOUT VOUT m1_9368_n744#
+ VDD VOUT m1_9368_n744# VOUT m1_9368_n744# m1_9368_n744# VOUT VDD m1_9368_n744# m1_9368_n744#
+ VDD VOUT VDD VOUT m1_9368_n744# m1_9368_n744# m1_9368_n744# sky130_fd_pr__pfet_g5v0d10v5_8UL4MK
Xsky130_fd_pr__cap_mim_m3_1_BHK9HY_0 m1_9368_n744# m1_9368_n744# m1_10706_1822# m1_10706_1822#
+ m1_10706_1822# m1_9368_n744# sky130_fd_pr__cap_mim_m3_1_BHK9HY
Xsky130_fd_pr__nfet_g5v0d10v5_7WHXCK_0 VOUT w_7736_n902# VSS VSS VSS VSS VSS VSS VBIAS
+ VSS VOUT VSS VOUT VSS VSS VOUT VOUT VBIAS VSS w_7736_n902# w_7736_n902# VSS VOUT
+ VSS VSS VSS VSS VOUT VBIAS VSS VOUT VOUT w_7736_n902# VSS w_7736_n902# VSS VOUT
+ VSS VSS VBIAS VBIAS VBIAS sky130_fd_pr__nfet_g5v0d10v5_7WHXCK
XXM10 VINN VINN m1_4902_n766# m1_4902_n766# m1_4902_n766# w_4240_n902# m1_4902_n766#
+ w_4240_n902# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902#
+ m1_4902_n766# VINN m1_4902_n766# w_4240_n902# m1_4902_n766# VINN VINN m1_4902_n766#
+ m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# w_4240_n902# VINN VINN m1_4902_n766#
+ w_4240_n902# w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902#
+ w_4240_n902# w_4240_n902# VINN VINN m1_4902_n766# VINN VINN m1_4902_n766# VINN VINN
+ m1_4902_n766# VINN m1_4902_n766# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN
+ VINN m1_4902_n766# w_4240_n902# m1_4902_n766# m1_4902_n766# m1_4902_n766# VINN m1_4902_n766#
+ VINN m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# m1_4902_n766# w_4240_n902#
+ VINN w_4240_n902# VINN w_4240_n902# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_KWU84Z a_n29_n2720# a_3067_1720# a_n287_610#
+ a_1261_n500# a_487_n1610# a_1777_1720# a_n2609_1720# a_n803_n2720# a_229_n2720#
+ a_n287_n1610# a_2867_n2808# a_n2351_1720# a_n1319_n500# a_n3125_610# a_n2609_610#
+ a_n287_n500# a_3067_n2720# a_229_1720# a_n1061_n500# a_n1577_1720# a_n3259_n2942#
+ a_2093_n2808# a_2551_610# a_2035_1720# a_n2351_n2720# a_1577_n2808# a_2551_n2720#
+ a_803_n2808# a_n745_n2808# a_n1003_n2808# a_3067_610# a_2809_n500# a_n1835_n2720#
+ a_745_n500# a_2035_610# a_n545_1720# a_1519_610# a_1003_610# a_745_n1610# a_2551_n500#
+ a_n1061_n2720# a_n545_n1610# a_1003_n1610# a_1261_n2720# a_3067_n500# a_1777_n500#
+ a_n2609_n500# a_1003_1720# a_n2293_n2808# a_n2867_n1610# a_n3125_n2720# a_n2351_610#
+ a_n2867_610# a_n1835_610# a_n2609_n2720# a_n1777_n2808# a_n2351_n500# a_2809_n2720#
+ a_2351_n2808# a_n2867_1720# a_n1319_610# a_1835_n2808# a_n803_610# a_229_n500# a_n2093_n1610#
+ a_2293_n1610# a_n1577_n500# a_n1577_n1610# a_2293_610# a_2035_n2720# a_n229_n2808#
+ a_1261_610# a_1777_610# a_2035_n500# a_n29_n1610# a_1777_n1610# a_n1319_n2720# a_n29_1720#
+ a_1519_n2720# a_487_1720# a_n3067_n2808# a_1061_n2808# a_n803_n1610# a_n545_n500#
+ a_229_n1610# a_487_n2720# a_2293_1720# a_n3125_1720# a_745_610# a_n1835_1720# a_n2551_n2808#
+ a_n287_n2720# a_2609_n2808# a_229_610# a_3067_n1610# a_n803_1720# a_n2093_610# a_1003_n500#
+ a_1519_1720# a_n1577_610# a_n2351_n1610# a_n1061_610# a_n2093_1720# a_2551_n1610#
+ a_n1261_n2808# a_n1835_n1610# a_1319_n2808# a_n2867_n500# a_1261_1720# a_n545_610#
+ a_287_n2808# a_n2809_n2808# a_745_n2720# a_n1061_n1610# a_n1319_1720# a_n29_n500#
+ a_1261_n1610# a_n545_n2720# a_487_n500# a_1003_n2720# a_n287_1720# a_n3125_n1610#
+ a_n1061_1720# a_487_610# a_n3125_n500# a_2293_n500# a_n2035_n2808# a_n2609_n1610#
+ a_n2867_n2720# a_n1835_n500# a_2809_n1610# a_n1519_n2808# a_2809_1720# a_n29_610#
+ a_745_1720# a_2809_610# a_n803_n500# a_n2093_n2720# a_2551_1720# a_1519_n500# a_2035_n1610#
+ a_545_n2808# a_n1319_n1610# a_2293_n2720# a_29_n2808# a_n487_n2808# a_n2093_n500#
+ a_n1577_n2720# a_1519_n1610# a_1777_n2720#
X0 a_n1061_1720# a_n1261_n2808# a_n1319_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X1 a_2551_n2720# a_2351_n2808# a_2293_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_1003_n500# a_803_n2808# a_745_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_n803_610# a_n1003_n2808# a_n1061_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a_n1835_n2720# a_n2035_n2808# a_n2093_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X5 a_n803_n1610# a_n1003_n2808# a_n1061_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X6 a_745_610# a_545_n2808# a_487_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X7 a_1003_1720# a_803_n2808# a_745_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X8 a_745_n500# a_545_n2808# a_487_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X9 a_n29_610# a_n229_n2808# a_n287_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X10 a_1261_n2720# a_1061_n2808# a_1003_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X11 a_745_1720# a_545_n2808# a_487_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X12 a_487_n500# a_287_n2808# a_229_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X13 a_487_1720# a_287_n2808# a_229_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X14 a_229_n2720# a_29_n2808# a_n29_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X15 a_n545_n2720# a_n745_n2808# a_n803_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X16 a_229_610# a_29_n2808# a_n29_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X17 a_2035_n500# a_1835_n2808# a_1777_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X18 a_3067_n1610# a_2867_n2808# a_2809_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X19 a_2035_1720# a_1835_n2808# a_1777_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X20 a_1777_n500# a_1577_n2808# a_1519_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X21 a_n2609_n500# a_n2809_n2808# a_n2867_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X22 a_1777_1720# a_1577_n2808# a_1519_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X23 a_n2609_1720# a_n2809_n2808# a_n2867_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X24 a_2809_n1610# a_2609_n2808# a_2551_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X25 a_1519_610# a_1319_n2808# a_1261_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X26 a_1777_n1610# a_1577_n2808# a_1519_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X27 a_1261_n500# a_1061_n2808# a_1003_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X28 a_1261_1720# a_1061_n2808# a_1003_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X29 a_n1835_n500# a_n2035_n2808# a_n2093_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X30 a_1519_n1610# a_1319_n2808# a_1261_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X31 a_487_610# a_287_n2808# a_229_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X32 a_n1835_1720# a_n2035_n2808# a_n2093_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X33 a_n2351_n2720# a_n2551_n2808# a_n2609_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X34 a_1003_n2720# a_803_n2808# a_745_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X35 a_2809_610# a_2609_n2808# a_2551_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X36 a_n545_610# a_n745_n2808# a_n803_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X37 a_n2867_n1610# a_n3067_n2808# a_n3125_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X38 a_n1061_n2720# a_n1261_n2808# a_n1319_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X39 a_n1319_610# a_n1519_n2808# a_n1577_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X40 a_487_n1610# a_287_n2808# a_229_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X41 a_2293_n1610# a_2093_n2808# a_2035_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X42 a_n1835_610# a_n2035_n2808# a_n2093_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X43 a_n803_n2720# a_n1003_n2808# a_n1061_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X44 a_1261_610# a_1061_n2808# a_1003_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X45 a_2809_n500# a_2609_n2808# a_2551_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X46 a_2809_1720# a_2609_n2808# a_2551_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X47 a_n287_n1610# a_n487_n2808# a_n545_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X48 a_n2609_610# a_n2809_n2808# a_n2867_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X49 a_n2351_n500# a_n2551_n2808# a_n2609_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X50 a_n2609_n1610# a_n2809_n2808# a_n2867_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X51 a_n2351_1720# a_n2551_n2808# a_n2609_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X52 a_n2093_n500# a_n2293_n2808# a_n2351_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X53 a_2035_610# a_1835_n2808# a_1777_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X54 a_n29_n1610# a_n229_n2808# a_n287_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X55 a_n1577_n1610# a_n1777_n2808# a_n1835_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X56 a_229_n500# a_29_n2808# a_n29_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X57 a_n2093_1720# a_n2293_n2808# a_n2351_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X58 a_n29_n500# a_n229_n2808# a_n287_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X59 a_229_1720# a_29_n2808# a_n29_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X60 a_3067_n2720# a_2867_n2808# a_2809_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X61 a_2035_n1610# a_1835_n2808# a_1777_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X62 a_2551_610# a_2351_n2808# a_2293_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X63 a_n29_1720# a_n229_n2808# a_n287_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X64 a_n1319_n1610# a_n1519_n2808# a_n1577_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X65 a_n1061_610# a_n1261_n2808# a_n1319_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X66 a_2809_n2720# a_2609_n2808# a_2551_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X67 a_n287_610# a_n487_n2808# a_n545_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X68 a_1777_n2720# a_1577_n2808# a_1519_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X69 a_1519_n2720# a_1319_n2808# a_1261_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X70 a_n2093_n1610# a_n2293_n2808# a_n2351_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X71 a_745_n1610# a_545_n2808# a_487_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X72 a_n2351_610# a_n2551_n2808# a_n2609_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X73 a_3067_n500# a_2867_n2808# a_2809_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X74 a_2551_n1610# a_2351_n2808# a_2293_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X75 a_3067_1720# a_2867_n2808# a_2809_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X76 a_n2867_n2720# a_n3067_n2808# a_n3125_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X77 a_n1835_n1610# a_n2035_n2808# a_n2093_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X78 a_487_n2720# a_287_n2808# a_229_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X79 a_2551_n500# a_2351_n2808# a_2293_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X80 a_n1319_n500# a_n1519_n2808# a_n1577_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X81 a_2293_n2720# a_2093_n2808# a_2035_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X82 a_1261_n1610# a_1061_n2808# a_1003_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X83 a_n2867_610# a_n3067_n2808# a_n3125_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X84 a_2293_n500# a_2093_n2808# a_2035_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X85 a_n545_n500# a_n745_n2808# a_n803_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X86 a_1777_610# a_1577_n2808# a_1519_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X87 a_n1319_1720# a_n1519_n2808# a_n1577_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X88 a_2551_1720# a_2351_n2808# a_2293_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X89 a_n287_n500# a_n487_n2808# a_n545_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X90 a_n545_1720# a_n745_n2808# a_n803_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X91 a_2293_1720# a_2093_n2808# a_2035_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X92 a_2293_610# a_2093_n2808# a_2035_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X93 a_229_n1610# a_29_n2808# a_n29_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X94 a_n545_n1610# a_n745_n2808# a_n803_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X95 a_n803_n500# a_n1003_n2808# a_n1061_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X96 a_n2867_n500# a_n3067_n2808# a_n3125_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X97 a_n287_1720# a_n487_n2808# a_n545_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X98 a_n2867_1720# a_n3067_n2808# a_n3125_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X99 a_n803_1720# a_n1003_n2808# a_n1061_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X100 a_n287_n2720# a_n487_n2808# a_n545_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X101 a_1003_610# a_803_n2808# a_745_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X102 a_n2609_n2720# a_n2809_n2808# a_n2867_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X103 a_3067_610# a_2867_n2808# a_2809_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X104 a_n29_n2720# a_n229_n2808# a_n287_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X105 a_n1577_n2720# a_n1777_n2808# a_n1835_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X106 a_n1577_610# a_n1777_n2808# a_n1835_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X107 a_2035_n2720# a_1835_n2808# a_1777_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X108 a_n2093_610# a_n2293_n2808# a_n2351_610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X109 a_n1319_n2720# a_n1519_n2808# a_n1577_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X110 a_n2351_n1610# a_n2551_n2808# a_n2609_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X111 a_n1577_n500# a_n1777_n2808# a_n1835_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X112 a_1003_n1610# a_803_n2808# a_745_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X113 a_1519_n500# a_1319_n2808# a_1261_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X114 a_n1577_1720# a_n1777_n2808# a_n1835_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X115 a_1519_1720# a_1319_n2808# a_1261_1720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X116 a_n2093_n2720# a_n2293_n2808# a_n2351_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X117 a_n1061_n1610# a_n1261_n2808# a_n1319_n1610# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X118 a_n1061_n500# a_n1261_n2808# a_n1319_n500# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X119 a_745_n2720# a_545_n2808# a_487_n2720# a_n3259_n2942# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt Input_Stage_OA2 VDD VOUT VINN VINP VBIAS w_8718_n902# w_7736_n902# VSS w_4240_n902#
XXR1 VSS m1_10706_1822# VOUT sky130_fd_pr__res_high_po_0p69_FJD3D2
Xsky130_fd_pr__nfet_05v0_nvt_FEJX3A_0 VINP VINP w_8718_n902# w_8718_n902# w_8718_n902#
+ m1_9368_n744# w_8718_n902# m1_9368_n744# w_8718_n902# VINP m1_9368_n744# m1_9368_n744#
+ VINP m1_9368_n744# m1_9368_n744# w_8718_n902# VINP w_8718_n902# m1_9368_n744# w_8718_n902#
+ VINP VINP w_8718_n902# w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902# w_8718_n902#
+ VINP VINP w_8718_n902# m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP m1_9368_n744#
+ m1_9368_n744# VINP m1_9368_n744# m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902#
+ VINP VINP w_8718_n902# VINP VINP w_8718_n902# VINP w_8718_n902# w_8718_n902# VINP
+ m1_9368_n744# m1_9368_n744# VINP VINP w_8718_n902# m1_9368_n744# w_8718_n902# w_8718_n902#
+ w_8718_n902# VINP w_8718_n902# VINP w_8718_n902# m1_9368_n744# m1_9368_n744# w_8718_n902#
+ w_8718_n902# m1_9368_n744# VINP m1_9368_n744# VINP m1_9368_n744# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
XXM2 VINN w_8718_n902# VINP w_7736_n902# w_7736_n902# w_4240_n902# w_7736_n902# sky130_fd_pr__nfet_01v8_lvt_AJ3MPE
XXM6 m1_9368_n744# m1_4902_n766# m1_9368_n744# VDD m1_4902_n766# m1_4902_n766# VDD
+ m1_4902_n766# m1_4902_n766# m1_4902_n766# VDD sky130_fd_pr__pfet_01v8_lvt_UX3DP3
XXM8 VDD VOUT VDD VOUT VDD VDD VOUT VDD m1_9368_n744# VDD VDD VOUT VOUT m1_9368_n744#
+ VDD VOUT m1_9368_n744# VOUT m1_9368_n744# m1_9368_n744# VOUT VDD m1_9368_n744# m1_9368_n744#
+ VDD VOUT VDD VOUT m1_9368_n744# m1_9368_n744# m1_9368_n744# sky130_fd_pr__pfet_g5v0d10v5_8UL4MK
Xsky130_fd_pr__cap_mim_m3_1_BHK9HY_0 m1_9368_n744# m1_9368_n744# m1_10706_1822# m1_10706_1822#
+ m1_10706_1822# m1_9368_n744# sky130_fd_pr__cap_mim_m3_1_BHK9HY
XXM10 VINN VINN m1_4902_n766# m1_4902_n766# m1_4902_n766# w_4240_n902# m1_4902_n766#
+ w_4240_n902# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902#
+ m1_4902_n766# VINN m1_4902_n766# w_4240_n902# m1_4902_n766# VINN VINN m1_4902_n766#
+ m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# w_4240_n902# VINN VINN m1_4902_n766#
+ w_4240_n902# w_4240_n902# w_4240_n902# VINN w_4240_n902# w_4240_n902# VINN w_4240_n902#
+ w_4240_n902# w_4240_n902# VINN VINN m1_4902_n766# VINN VINN m1_4902_n766# VINN VINN
+ m1_4902_n766# VINN m1_4902_n766# m1_4902_n766# VINN w_4240_n902# w_4240_n902# VINN
+ VINN m1_4902_n766# w_4240_n902# m1_4902_n766# m1_4902_n766# m1_4902_n766# VINN m1_4902_n766#
+ VINN m1_4902_n766# w_4240_n902# w_4240_n902# m1_4902_n766# m1_4902_n766# w_4240_n902#
+ VINN w_4240_n902# VINN w_4240_n902# sky130_fd_pr__nfet_05v0_nvt_FEJX3A
Xsky130_fd_pr__nfet_g5v0d10v5_KWU84Z_0 VSS VSS VOUT VOUT VSS VOUT VSS VOUT VOUT VOUT
+ VBIAS VOUT VOUT VSS VSS VOUT VSS VOUT VSS VSS VSS VBIAS VSS VSS VOUT VBIAS VSS VBIAS
+ VBIAS VBIAS VSS w_7736_n902# VOUT VOUT VSS VSS VSS VSS VOUT VSS VSS VSS VSS VOUT
+ VSS VOUT VSS VSS VBIAS VOUT VSS VOUT VOUT VOUT VSS VBIAS VOUT w_7736_n902# VBIAS
+ VOUT VOUT VBIAS VOUT VOUT VSS w_7736_n902# VSS VSS w_7736_n902# VSS VBIAS VOUT VOUT
+ VSS VSS VOUT VOUT VSS VSS VSS VBIAS VBIAS VOUT VSS VOUT VSS w_7736_n902# VSS VOUT
+ VOUT VBIAS VOUT VBIAS VOUT VSS VOUT VSS VSS VSS VSS VOUT VSS VSS VSS VBIAS VOUT
+ VBIAS VOUT VOUT VSS VBIAS VBIAS VOUT VSS VOUT VSS VOUT VSS VSS VSS VOUT VSS VSS
+ VSS VSS w_7736_n902# VBIAS VSS VOUT VOUT w_7736_n902# VBIAS w_7736_n902# VSS VOUT
+ w_7736_n902# VOUT VSS VSS VSS VSS VBIAS VOUT w_7736_n902# VBIAS VBIAS VSS VSS VSS
+ VOUT sky130_fd_pr__nfet_g5v0d10v5_KWU84Z
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_TVN32V a_3368_n2141# a_n118_1709# a_48_n2141#
+ a_n2774_1709# a_1542_1709# a_n2940_n2141# a_n782_1709# a_2372_n2141# a_3700_n2141#
+ a_n1944_n2141# a_n3106_1709# a_n3438_n2141# a_n782_n2141# a_n1280_1709# a_1376_1709#
+ a_1376_n2141# a_2704_n2141# a_546_n2141# a_n2608_1709# a_380_1709# a_n3770_1709#
+ a_1708_n2141# a_3866_1709# a_n2442_n2141# a_n616_1709# a_4198_1709# a_3202_n2141#
+ a_n1446_n2141# a_n1114_1709# a_n4102_1709# a_n284_n2141# a_2206_n2141# a_2372_1709#
+ a_214_1709# a_n3604_1709# a_n616_n2141# a_1874_1709# a_1210_n2141# a_n3438_1709#
+ a_n2110_1709# a_2206_1709# a_4198_n2141# a_48_1709# a_878_n2141# a_n118_n2141# a_n1612_1709#
+ a_n3770_n2141# a_1708_1709# a_2870_1709# a_712_1709# a_n2774_n2141# a_n948_1709#
+ a_n4268_n2141# a_3534_n2141# a_n1778_n2141# a_n1446_1709# a_3202_1709# a_2538_n2141#
+ a_546_1709# a_n3272_n2141# a_n3936_1709# a_n948_n2141# a_2704_1709# a_380_n2141#
+ a_4032_n2141# a_n2276_n2141# a_n3604_n2141# a_n4268_1709# a_1542_n2141# a_3036_1709#
+ a_712_n2141# a_3036_n2141# a_n2608_n2141# a_n2442_1709# a_2538_1709# a_1210_1709#
+ a_n1280_n2141# a_n4102_n2141# a_n1944_1709# a_n450_1709# a_2040_n2141# a_3700_1709#
+ a_n1612_n2141# a_n450_n2141# a_n2276_1709# a_n3106_n2141# a_1044_1709# a_1044_n2141#
+ a_4032_1709# a_214_n2141# a_3866_n2141# a_n1778_1709# a_n284_1709# a_3534_1709#
+ a_n4398_n2271# a_n2110_n2141# a_878_1709# a_n2940_1709# a_n1114_n2141# a_2870_n2141#
+ a_n3272_1709# a_n3936_n2141# a_1874_n2141# a_2040_1709# a_3368_1709#
X0 a_n782_1709# a_n782_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X1 a_1376_1709# a_1376_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X2 a_4198_1709# a_4198_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X3 a_878_1709# a_878_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X4 a_n3770_1709# a_n3770_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X5 a_n1446_1709# a_n1446_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X6 a_3700_1709# a_3700_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X7 a_n4268_1709# a_n4268_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X8 a_n2110_1709# a_n2110_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X9 a_1874_1709# a_1874_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X10 a_2372_1709# a_2372_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X11 a_2538_1709# a_2538_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X12 a_3036_1709# a_3036_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X13 a_n1944_1709# a_n1944_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X14 a_214_1709# a_214_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X15 a_n2608_1709# a_n2608_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X16 a_n2442_1709# a_n2442_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X17 a_n3106_1709# a_n3106_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X18 a_2870_1709# a_2870_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X19 a_1210_1709# a_1210_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X20 a_3534_1709# a_3534_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X21 a_n1280_1709# a_n1280_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X22 a_4032_1709# a_4032_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X23 a_712_1709# a_712_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X24 a_n3604_1709# a_n3604_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X25 a_n118_1709# a_n118_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X26 a_n4102_1709# a_n4102_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X27 a_n1778_1709# a_n1778_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X28 a_n2276_1709# a_n2276_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X29 a_n616_1709# a_n616_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X30 a_1044_1709# a_1044_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X31 a_3368_1709# a_3368_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X32 a_380_1709# a_380_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X33 a_546_1709# a_546_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X34 a_n2940_1709# a_n2940_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X35 a_n2774_1709# a_n2774_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X36 a_n3438_1709# a_n3438_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X37 a_n3272_1709# a_n3272_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X38 a_n1114_1709# a_n1114_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X39 a_1542_1709# a_1542_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X40 a_1708_1709# a_1708_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X41 a_3866_1709# a_3866_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X42 a_2040_1709# a_2040_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X43 a_2206_1709# a_2206_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X44 a_n3936_1709# a_n3936_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X45 a_n1612_1709# a_n1612_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X46 a_n450_1709# a_n450_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X47 a_n284_1709# a_n284_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X48 a_48_1709# a_48_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X49 a_2704_1709# a_2704_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X50 a_n948_1709# a_n948_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
X51 a_3202_1709# a_3202_n2141# a_n4398_n2271# sky130_fd_pr__res_xhigh_po_0p35 l=17.25
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_QHQRGL a_1044_n2396# a_214_n2396# a_n1446_1964#
+ a_546_1964# a_n2110_n2396# a_n1114_n2396# a_n2406_n2526# a_1874_n2396# a_1210_1964#
+ a_48_n2396# a_n1944_1964# a_n450_1964# a_1044_1964# a_n1944_n2396# a_n2276_1964#
+ a_1376_n2396# a_n782_n2396# a_n1778_1964# a_546_n2396# a_n284_1964# a_1708_n2396#
+ a_878_1964# a_2040_1964# a_n1446_n2396# a_2206_n2396# a_n118_1964# a_n284_n2396#
+ a_1542_1964# a_n616_n2396# a_n782_1964# a_1210_n2396# a_1376_1964# a_n1280_1964#
+ a_380_1964# a_878_n2396# a_n118_n2396# a_n616_1964# a_n1114_1964# a_214_1964# a_n1778_n2396#
+ a_1874_1964# a_n948_n2396# a_380_n2396# a_n2276_n2396# a_2206_1964# a_1542_n2396#
+ a_712_n2396# a_n2110_1964# a_48_1964# a_1708_1964# a_n1280_n2396# a_n1612_1964#
+ a_2040_n2396# a_712_1964# a_n1612_n2396# a_n450_n2396# a_n948_1964#
X0 a_1874_1964# a_1874_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X1 a_n1944_1964# a_n1944_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X2 a_214_1964# a_214_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X3 a_1210_1964# a_1210_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X4 a_n1280_1964# a_n1280_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X5 a_712_1964# a_712_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X6 a_n118_1964# a_n118_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X7 a_n1778_1964# a_n1778_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X8 a_n2276_1964# a_n2276_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X9 a_n616_1964# a_n616_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X10 a_1044_1964# a_1044_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X11 a_380_1964# a_380_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X12 a_546_1964# a_546_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X13 a_n1114_1964# a_n1114_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X14 a_1542_1964# a_1542_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X15 a_1708_1964# a_1708_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X16 a_2040_1964# a_2040_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X17 a_2206_1964# a_2206_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X18 a_n1612_1964# a_n1612_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X19 a_n450_1964# a_n450_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X20 a_n284_1964# a_n284_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X21 a_48_1964# a_48_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X22 a_n948_1964# a_n948_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X23 a_n782_1964# a_n782_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X24 a_1376_1964# a_1376_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X25 a_878_1964# a_878_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X26 a_n1446_1964# a_n1446_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
X27 a_n2110_1964# a_n2110_n2396# a_n2406_n2526# sky130_fd_pr__res_xhigh_po_0p35 l=19.8
.ends

.subckt Input_Stage_v1 VINP VOUT1 VINN CM VBIAS w_18276_n26882# w_22762_n17134# w_21780_n17134#
+ w_21772_n36602# w_22754_n36602# w_18284_n17134# w_21772_n26882# w_22754_n26882#
+ w_18276_n36602# AVDD AVSS
Xx1 AVDD x1/VOUT x1/VOUT VINN VBIAS w_22754_n36602# w_21772_n36602# AVSS w_18276_n36602#
+ Input_Stage_OA1
Xx2 AVDD x2/VOUT x2/VOUT VINP VBIAS w_22754_n26882# w_21772_n26882# AVSS w_18276_n26882#
+ Input_Stage_OA1
Xx3 AVDD VOUT1 x3/VINN x3/VINP VBIAS w_22762_n17134# w_21780_n17134# AVSS w_18284_n17134#
+ Input_Stage_OA2
Xsky130_fd_pr__res_xhigh_po_0p35_TVN32V_0 m1_23074_n22690# m1_19588_n18840# m1_19754_n22690#
+ m1_16932_n18840# m1_21248_n18840# m1_16766_n22690# m1_18924_n18840# m1_22078_n22690#
+ m1_23406_n22690# m1_17762_n22690# m1_16600_n18840# m1_16434_n22690# m1_19090_n22690#
+ m1_18592_n18840# m1_21248_n18840# m1_21082_n22690# m1_22410_n22690# m1_20418_n22690#
+ m1_17264_n18840# m1_20252_n18840# m1_15936_n18840# m1_21414_n22690# m1_23572_n18840#
+ m1_17430_n22690# m1_19256_n18840# m1_23904_n18840# m1_23074_n22690# m1_18426_n22690#
+ m1_18592_n18840# x3/VINP m1_19422_n22690# m1_22078_n22690# m1_22244_n18840# m1_19920_n18840#
+ m1_16268_n18840# m1_19090_n22690# m1_21580_n18840# m1_21082_n22690# m1_16268_n18840#
+ m1_17596_n18840# m1_21912_n18840# VINP m1_19920_n18840# m1_20750_n22690# m1_19754_n22690#
+ m1_18260_n18840# m1_16102_n22690# m1_21580_n18840# m1_22576_n18840# m1_20584_n18840#
+ m1_17098_n22690# m1_18924_n18840# m1_15606_n22692# m1_23406_n22690# m1_18094_n22690#
+ m1_18260_n18840# m1_22908_n18840# m1_22410_n22690# m1_20252_n18840# m1_16434_n22690#
+ m1_15936_n18840# m1_18758_n22690# m1_22576_n18840# m1_20086_n22690# m1_23738_n22690#
+ m1_17430_n22690# m1_16102_n22690# x2/VOUT m1_21414_n22690# m1_22908_n18840# m1_20418_n22690#
+ m1_22742_n22690# m1_17098_n22690# m1_17264_n18840# m1_22244_n18840# m1_20916_n18840#
+ m1_18426_n22690# m1_15606_n22692# m1_17928_n18840# m1_19256_n18840# m1_21746_n22690#
+ m1_23572_n18840# m1_18094_n22690# m1_19422_n22690# m1_17596_n18840# m1_16766_n22690#
+ m1_20916_n18840# m1_20750_n22690# m1_23904_n18840# m1_20086_n22690# m1_23738_n22690#
+ m1_17928_n18840# m1_19588_n18840# m1_23240_n18840# AVSS m1_17762_n22690# m1_20584_n18840#
+ m1_16932_n18840# m1_18758_n22690# m1_22742_n22690# m1_16600_n18840# CM m1_21746_n22690#
+ m1_21912_n18840# m1_23240_n18840# sky130_fd_pr__res_xhigh_po_0p35_TVN32V
Xsky130_fd_pr__res_xhigh_po_0p35_TVN32V_1 m1_23104_n32408# m1_19618_n28558# m1_19784_n32408#
+ m1_16962_n28558# m1_21278_n28558# m1_16796_n32408# m1_18954_n28558# m1_22108_n32408#
+ m1_23436_n32408# m1_17792_n32408# m1_16630_n28558# m1_16464_n32408# m1_19120_n32408#
+ m1_18622_n28558# m1_21278_n28558# m1_21112_n32408# m1_22440_n32408# m1_20448_n32408#
+ m1_17294_n28558# m1_20282_n28558# m1_15966_n28558# m1_21444_n32408# m1_23602_n28558#
+ m1_17460_n32408# m1_19286_n28558# m1_23934_n28558# m1_23104_n32408# m1_18456_n32408#
+ m1_18622_n28558# x3/VINN m1_19452_n32408# m1_22108_n32408# m1_22274_n28558# m1_19950_n28558#
+ m1_16298_n28558# m1_19120_n32408# m1_21610_n28558# m1_21112_n32408# m1_16298_n28558#
+ m1_17626_n28558# m1_21942_n28558# VINN m1_19950_n28558# m1_20780_n32408# m1_19784_n32408#
+ m1_18290_n28558# m1_16132_n32408# m1_21610_n28558# m1_22606_n28558# m1_20614_n28558#
+ m1_17128_n32408# m1_18954_n28558# m1_15634_n32408# m1_23436_n32408# m1_18124_n32408#
+ m1_18290_n28558# m1_22938_n28558# m1_22440_n32408# m1_20282_n28558# m1_16464_n32408#
+ m1_15966_n28558# m1_18788_n32408# m1_22606_n28558# m1_20116_n32408# m1_23768_n32408#
+ m1_17460_n32408# m1_16132_n32408# x1/VOUT m1_21444_n32408# m1_22938_n28558# m1_20448_n32408#
+ m1_22772_n32408# m1_17128_n32408# m1_17294_n28558# m1_22274_n28558# m1_20946_n28558#
+ m1_18456_n32408# m1_15634_n32408# m1_17958_n28558# m1_19286_n28558# m1_21776_n32408#
+ m1_23602_n28558# m1_18124_n32408# m1_19452_n32408# m1_17626_n28558# m1_16796_n32408#
+ m1_20946_n28558# m1_20780_n32408# m1_23934_n28558# m1_20116_n32408# m1_23768_n32408#
+ m1_17958_n28558# m1_19618_n28558# m1_23270_n28558# AVSS m1_17792_n32408# m1_20614_n28558#
+ m1_16962_n28558# m1_18788_n32408# m1_22772_n32408# m1_16630_n28558# CM m1_21776_n32408#
+ m1_21942_n28558# m1_23270_n28558# sky130_fd_pr__res_xhigh_po_0p35_TVN32V
Xsky130_fd_pr__res_xhigh_po_0p35_QHQRGL_0 m1_18184_n12946# m1_17520_n12946# m1_15694_n8586#
+ m1_17686_n8586# m1_15196_n12946# m1_16192_n12946# AVSS m1_19180_n12946# m1_18350_n8586#
+ CM m1_15362_n8586# m1_16690_n8586# m1_18350_n8586# m1_15196_n12946# m1_15030_n8586#
+ m1_18516_n12946# m1_16524_n12946# m1_15362_n8586# m1_17852_n12946# m1_17022_n8586#
+ m1_18848_n12946# m1_18018_n8586# m1_19346_n8586# m1_15860_n12946# x3/VINP m1_17022_n8586#
+ m1_16856_n12946# m1_18682_n8586# m1_16524_n12946# m1_16358_n8586# m1_18516_n12946#
+ m1_18682_n8586# m1_16026_n8586# m1_17686_n8586# m1_18184_n12946# x3/VINN m1_16690_n8586#
+ m1_16026_n8586# m1_17354_n8586# m1_15528_n12946# m1_19014_n8586# m1_16192_n12946#
+ m1_17520_n12946# VOUT1 m1_19346_n8586# m1_18848_n12946# m1_17852_n12946# m1_15030_n8586#
+ m1_17354_n8586# m1_19014_n8586# m1_15860_n12946# m1_15694_n8586# m1_19180_n12946#
+ m1_18018_n8586# m1_15528_n12946# m1_16856_n12946# m1_16358_n8586# sky130_fd_pr__res_xhigh_po_0p35_QHQRGL
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TZT4V2 a_100_n500# a_n292_n722# a_n158_n500#
+ a_n100_n588#
X0 a_100_n500# a_n100_n588# a_n158_n500# a_n292_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
.ends

.subckt vbias_gen_pga VBIAS IBIAS VSS
XXM4 VSS VSS VBIAS VBIAS sky130_fd_pr__nfet_g5v0d10v5_TZT4V2
R0 IBIAS VBIAS sky130_fd_pr__res_generic_m1 w=1 l=0.08
.ends

.subckt sky130_pa_ip__instramp V[9] V[8] V[7] V[6] V[5] V[4] V[3] V[2] V[1] V[0] VCM
+ IBIAS VINP DVDD VOUT VINN w_6926_14586# w_3442_14586# w_21944_24334# w_7900_24334#
+ w_3442_4866# w_21946_14614# w_7908_14586# w_22926_24334# w_18448_24334# w_7908_4866#
+ w_21948_4866# w_6918_24334# w_3434_24334# w_22928_14614# w_22930_4866# w_18452_4866#
+ w_18450_14614# w_6926_4866# AVDD AVSS DVSS
Xx1 V[6] V[5] V[8] V[9] V[7] x1/VO1 VOUT V[4] V[3] V[2] V[1] V[0] VCM w_18452_4866#
+ x3/VBIAS w_18448_24334# w_22928_14614# w_22930_4866# w_18450_14614# w_22926_24334#
+ DVDD w_21948_4866# w_21946_14614# DVSS AVSS AVDD w_21944_24334# Parallel_10B_Block2
Xx2 VINP x1/VO1 VINN VCM x3/VBIAS w_7908_14586# w_3434_24334# w_6918_24334# w_6926_4866#
+ w_3442_4866# w_7900_24334# w_6926_14586# w_3442_14586# w_7908_4866# AVDD AVSS Input_Stage_v1
Xx3 x3/VBIAS IBIAS AVSS vbias_gen_pga
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_N9BQ2J a_n345_n500# a_129_n500# a_287_n500# a_n479_n722#
+ a_29_n588# a_n129_n588# a_187_n588# a_n287_n588# a_n29_n500# a_n187_n500#
X0 a_n187_n500# a_n287_n588# a_n345_n500# a_n479_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X1 a_287_n500# a_187_n588# a_129_n500# a_n479_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X2 a_129_n500# a_29_n588# a_n29_n500# a_n479_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X3 a_n29_n500# a_n129_n588# a_n187_n500# a_n479_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLJ6Y6 a_n345_n500# a_29_n597# a_n129_n597# a_187_n597#
+ a_n503_n500# a_129_n500# a_n287_n597# w_n861_n797# a_287_n500# a_n661_n500# a_345_n597#
+ a_n445_n597# a_445_n500# a_503_n597# a_n603_n597# a_603_n500# a_n29_n500# a_n187_n500#
X0 a_n187_n500# a_n287_n597# a_n345_n500# w_n861_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X1 a_287_n500# a_187_n597# a_129_n500# w_n861_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X2 a_n345_n500# a_n445_n597# a_n503_n500# w_n861_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X3 a_129_n500# a_29_n597# a_n29_n500# w_n861_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X4 a_445_n500# a_345_n597# a_287_n500# w_n861_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X5 a_n503_n500# a_n603_n597# a_n661_n500# w_n861_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X6 a_n29_n500# a_n129_n597# a_n187_n500# w_n861_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X7 a_603_n500# a_503_n597# a_445_n500# w_n861_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
.ends

.subckt simple_analog_switch_2 on vdd vss off out in
XXM15 in out in vss on on on on in out sky130_fd_pr__nfet_g5v0d10v5_N9BQ2J
XXM4 out off off off in in off vdd out out off off in off off out out in sky130_fd_pr__pfet_g5v0d10v5_KLJ6Y6
.ends

.subckt sky130_fd_sc_hvl__inv_2 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X2 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X3 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt sky130_fd_sc_hvl__decap_4 VGND VNB VPB VPWR
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0 ps=0 w=0.75 l=1
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0 ps=0 w=1 l=1
.ends

.subckt simplest_analog_switch_ena1v8 avdd dvdd avss on out dvss in
Xsimple_analog_switch_2_0 sky130_fd_sc_hvl__inv_2_0/Y avdd avss sky130_fd_sc_hvl__inv_2_1/Y
+ out in simple_analog_switch_2
Xsky130_fd_sc_hvl__inv_2_0 sky130_fd_sc_hvl__inv_2_1/Y dvss dvss avdd avdd sky130_fd_sc_hvl__inv_2_0/Y
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_1 sky130_fd_sc_hvl__inv_2_1/A dvss dvss avdd avdd sky130_fd_sc_hvl__inv_2_1/Y
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 on dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_1/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__diode_2_0 on dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_0 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__decap_4_1 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
.ends

.subckt simple_switch_array_53 simplest_analog_switch_ena1v8_1[1]/on simplest_analog_switch_ena1v8_0[18]/on
+ simplest_analog_switch_ena1v8_0[27]/on simplest_analog_switch_ena1v8_2[1]/on simplest_analog_switch_ena1v8_2[2]/avdd
+ simplest_analog_switch_ena1v8_1[1]/dvdd simplest_analog_switch_ena1v8_3[1]/on simplest_analog_switch_ena1v8_2[0]/dvdd
+ simplest_analog_switch_ena1v8_0[15]/on simplest_analog_switch_ena1v8_0[24]/on simplest_analog_switch_ena1v8_6[1]/avdd
+ simplest_analog_switch_ena1v8_4[1]/on simplest_analog_switch_ena1v8_0[8]/on simplest_analog_switch_ena1v8_6[2]/avdd
+ simplest_analog_switch_ena1v8_1[0]/dvdd simplest_analog_switch_ena1v8_0[9]/avdd
+ simplest_analog_switch_ena1v8_5[1]/on simplest_analog_switch_ena1v8_0[26]/dvdd simplest_analog_switch_ena1v8_0[4]/avdd
+ simplest_analog_switch_ena1v8_0[12]/on simplest_analog_switch_ena1v8_0[21]/on simplest_analog_switch_ena1v8_2[1]/dvdd
+ simplest_analog_switch_ena1v8_3[0]/dvdd simplest_analog_switch_ena1v8_6[1]/on simplest_analog_switch_ena1v8_4[1]/dvdd
+ simplest_analog_switch_ena1v8_0[5]/on simplest_analog_switch_ena1v8_5[2]/dvdd simplest_analog_switch_ena1v8_7[1]/on
+ simplest_analog_switch_ena1v8_3[3]/avdd simplest_analog_switch_ena1v8_4[1]/avdd
+ simplest_analog_switch_ena1v8_7[1]/in simplest_analog_switch_ena1v8_2[3]/avdd simplest_analog_switch_ena1v8_0[2]/on
+ simplest_analog_switch_ena1v8_4[0]/dvdd simplest_analog_switch_ena1v8_1[2]/on simplest_analog_switch_ena1v8_0[19]/on
+ simplest_analog_switch_ena1v8_0[28]/on simplest_analog_switch_ena1v8_2[1]/in simplest_analog_switch_ena1v8_6[2]/dvdd
+ simplest_analog_switch_ena1v8_3[1]/dvdd simplest_analog_switch_ena1v8_2[2]/on simplest_analog_switch_ena1v8_5[3]/dvdd
+ simplest_analog_switch_ena1v8_4[0]/avdd simplest_analog_switch_ena1v8_0[4]/dvdd
+ simplest_analog_switch_ena1v8_5[2]/avdd simplest_analog_switch_ena1v8_3[2]/on simplest_analog_switch_ena1v8_0[25]/on
+ simplest_analog_switch_ena1v8_0[16]/on simplest_analog_switch_ena1v8_1[3]/dvdd simplest_analog_switch_ena1v8_1[3]/avdd
+ simplest_analog_switch_ena1v8_0[9]/on simplest_analog_switch_ena1v8_5[2]/on simplest_analog_switch_ena1v8_6[1]/in
+ simplest_analog_switch_ena1v8_7[0]/dvdd simplest_analog_switch_ena1v8_3[1]/avss
+ simplest_analog_switch_ena1v8_5[1]/avdd simplest_analog_switch_ena1v8_1[2]/dvdd
+ simplest_analog_switch_ena1v8_0[13]/on simplest_analog_switch_ena1v8_0[22]/on simplest_analog_switch_ena1v8_2[2]/dvdd
+ simplest_analog_switch_ena1v8_6[0]/dvdd simplest_analog_switch_ena1v8_2[3]/in simplest_analog_switch_ena1v8_6[2]/on
+ simplest_analog_switch_ena1v8_3[2]/dvdd simplest_analog_switch_ena1v8_1[1]/avdd
+ simplest_analog_switch_ena1v8_0[6]/on simplest_analog_switch_ena1v8_0[26]/avss simplest_analog_switch_ena1v8_2[0]/in
+ simplest_analog_switch_ena1v8_0[10]/on simplest_analog_switch_ena1v8_4[1]/out simplest_analog_switch_ena1v8_5[0]/in
+ simplest_analog_switch_ena1v8_0[3]/on simplest_analog_switch_ena1v8_0[29]/dvdd simplest_analog_switch_ena1v8_0[23]/avdd
+ simplest_analog_switch_ena1v8_1[0]/avdd simplest_analog_switch_ena1v8_5[1]/avss
+ simplest_analog_switch_ena1v8_0[2]/in simplest_analog_switch_ena1v8_2[0]/avdd simplest_analog_switch_ena1v8_2[3]/avss
+ simplest_analog_switch_ena1v8_1[3]/on simplest_analog_switch_ena1v8_0[29]/on simplest_analog_switch_ena1v8_4[0]/in
+ simplest_analog_switch_ena1v8_2[3]/on simplest_analog_switch_ena1v8_0[0]/on simplest_analog_switch_ena1v8_4[0]/avss
+ simplest_analog_switch_ena1v8_3[3]/on simplest_analog_switch_ena1v8_7[0]/in simplest_analog_switch_ena1v8_1[0]/on
+ simplest_analog_switch_ena1v8_0[19]/dvdd simplest_analog_switch_ena1v8_0[17]/on
+ simplest_analog_switch_ena1v8_0[26]/on simplest_analog_switch_ena1v8_0[23]/avss
+ simplest_analog_switch_ena1v8_0[14]/dvdd simplest_analog_switch_ena1v8_5[2]/avss
+ simplest_analog_switch_ena1v8_0[29]/avdd simplest_analog_switch_ena1v8_2[0]/on simplest_analog_switch_ena1v8_0[19]/avdd
+ simplest_analog_switch_ena1v8_5[0]/dvdd simplest_analog_switch_ena1v8_1[2]/avdd
+ simplest_analog_switch_ena1v8_0[9]/dvdd simplest_analog_switch_ena1v8_2[3]/out simplest_analog_switch_ena1v8_0[4]/avss
+ simplest_analog_switch_ena1v8_7[0]/avdd simplest_analog_switch_ena1v8_5[1]/dvdd
+ simplest_analog_switch_ena1v8_3[3]/avss simplest_analog_switch_ena1v8_3[2]/avdd
+ simplest_analog_switch_ena1v8_5[3]/on simplest_analog_switch_ena1v8_0[7]/in simplest_analog_switch_ena1v8_3[0]/on
+ simplest_analog_switch_ena1v8_0[14]/on simplest_analog_switch_ena1v8_3[0]/avdd simplest_analog_switch_ena1v8_0[23]/on
+ simplest_analog_switch_ena1v8_2[3]/dvdd simplest_analog_switch_ena1v8_3[3]/dvdd
+ simplest_analog_switch_ena1v8_4[1]/avss simplest_analog_switch_ena1v8_4[0]/on simplest_analog_switch_ena1v8_0[7]/on
+ simplest_analog_switch_ena1v8_1[0]/avss simplest_analog_switch_ena1v8_3[3]/out simplest_analog_switch_ena1v8_0[9]/avss
+ simplest_analog_switch_ena1v8_0[1]/in simplest_analog_switch_ena1v8_7[0]/avss simplest_analog_switch_ena1v8_1[2]/avss
+ simplest_analog_switch_ena1v8_7[1]/out simplest_analog_switch_ena1v8_5[3]/avdd simplest_analog_switch_ena1v8_5[0]/on
+ simplest_analog_switch_ena1v8_0[0]/in simplest_analog_switch_ena1v8_2[0]/avss simplest_analog_switch_ena1v8_3[2]/avss
+ simplest_analog_switch_ena1v8_1[3]/avss simplest_analog_switch_ena1v8_6[2]/avss
+ simplest_analog_switch_ena1v8_0[26]/avdd simplest_analog_switch_ena1v8_0[8]/in simplest_analog_switch_ena1v8_0[11]/on
+ simplest_analog_switch_ena1v8_3[1]/avdd simplest_analog_switch_ena1v8_0[20]/on simplest_analog_switch_ena1v8_2[1]/avdd
+ simplest_analog_switch_ena1v8_5[3]/out simplest_analog_switch_ena1v8_6[0]/on simplest_analog_switch_ena1v8_6[2]/in
+ simplest_analog_switch_ena1v8_0[23]/dvdd simplest_analog_switch_ena1v8_0[4]/on simplest_analog_switch_ena1v8_1[3]/out
+ simplest_analog_switch_ena1v8_6[1]/avss simplest_analog_switch_ena1v8_6[0]/in simplest_analog_switch_ena1v8_7[0]/on
+ simplest_analog_switch_ena1v8_3[0]/avss simplest_analog_switch_ena1v8_7[1]/dvdd
+ simplest_analog_switch_ena1v8_0[14]/avdd simplest_analog_switch_ena1v8_0[5]/in simplest_analog_switch_ena1v8_5[2]/in
+ simplest_analog_switch_ena1v8_0[29]/avss simplest_analog_switch_ena1v8_6[2]/out
+ simplest_analog_switch_ena1v8_6[0]/avss simplest_analog_switch_ena1v8_1[1]/avss
+ simplest_analog_switch_ena1v8_2[2]/avss simplest_analog_switch_ena1v8_6[0]/avdd
+ simplest_analog_switch_ena1v8_2[1]/avss simplest_analog_switch_ena1v8_7[1]/avdd
+ simplest_analog_switch_ena1v8_7[1]/avss simplest_analog_switch_ena1v8_5[0]/avss
+ simplest_analog_switch_ena1v8_0[14]/avss simplest_analog_switch_ena1v8_5[0]/avdd
+ simplest_analog_switch_ena1v8_0[1]/on simplest_analog_switch_ena1v8_0[19]/avss simplest_analog_switch_ena1v8_0[6]/in
+ simplest_analog_switch_ena1v8_5[3]/avss simplest_analog_switch_ena1v8_6[1]/dvdd
+ VSUBS
Xsimplest_analog_switch_ena1v8_0[0] simplest_analog_switch_ena1v8_2[0]/avdd simplest_analog_switch_ena1v8_2[0]/dvdd
+ simplest_analog_switch_ena1v8_2[0]/avss simplest_analog_switch_ena1v8_0[0]/on simplest_analog_switch_ena1v8_2[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[1] simplest_analog_switch_ena1v8_2[1]/avdd simplest_analog_switch_ena1v8_2[1]/dvdd
+ simplest_analog_switch_ena1v8_2[1]/avss simplest_analog_switch_ena1v8_0[1]/on simplest_analog_switch_ena1v8_2[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[2] simplest_analog_switch_ena1v8_2[2]/avdd simplest_analog_switch_ena1v8_2[2]/dvdd
+ simplest_analog_switch_ena1v8_2[2]/avss simplest_analog_switch_ena1v8_0[2]/on simplest_analog_switch_ena1v8_2[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[2]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[3] simplest_analog_switch_ena1v8_2[3]/avdd simplest_analog_switch_ena1v8_2[3]/dvdd
+ simplest_analog_switch_ena1v8_2[3]/avss simplest_analog_switch_ena1v8_0[3]/on simplest_analog_switch_ena1v8_2[3]/out
+ VSUBS simplest_analog_switch_ena1v8_6[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[4] simplest_analog_switch_ena1v8_0[4]/avdd simplest_analog_switch_ena1v8_0[4]/dvdd
+ simplest_analog_switch_ena1v8_0[4]/avss simplest_analog_switch_ena1v8_0[4]/on simplest_analog_switch_ena1v8_2[3]/out
+ VSUBS simplest_analog_switch_ena1v8_6[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[5] simplest_analog_switch_ena1v8_3[0]/avdd simplest_analog_switch_ena1v8_3[0]/dvdd
+ simplest_analog_switch_ena1v8_3[0]/avss simplest_analog_switch_ena1v8_0[5]/on simplest_analog_switch_ena1v8_3[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[5]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[6] simplest_analog_switch_ena1v8_3[1]/avdd simplest_analog_switch_ena1v8_3[1]/dvdd
+ simplest_analog_switch_ena1v8_3[1]/avss simplest_analog_switch_ena1v8_0[6]/on simplest_analog_switch_ena1v8_3[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[6]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[7] simplest_analog_switch_ena1v8_3[2]/avdd simplest_analog_switch_ena1v8_3[2]/dvdd
+ simplest_analog_switch_ena1v8_3[2]/avss simplest_analog_switch_ena1v8_0[7]/on simplest_analog_switch_ena1v8_3[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[7]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[8] simplest_analog_switch_ena1v8_3[3]/avdd simplest_analog_switch_ena1v8_3[3]/dvdd
+ simplest_analog_switch_ena1v8_3[3]/avss simplest_analog_switch_ena1v8_0[8]/on simplest_analog_switch_ena1v8_3[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[8]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[9] simplest_analog_switch_ena1v8_0[9]/avdd simplest_analog_switch_ena1v8_0[9]/dvdd
+ simplest_analog_switch_ena1v8_0[9]/avss simplest_analog_switch_ena1v8_0[9]/on simplest_analog_switch_ena1v8_3[3]/out
+ VSUBS simplest_analog_switch_ena1v8_4[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[10] simplest_analog_switch_ena1v8_1[0]/avdd simplest_analog_switch_ena1v8_1[0]/dvdd
+ simplest_analog_switch_ena1v8_1[0]/avss simplest_analog_switch_ena1v8_0[10]/on simplest_analog_switch_ena1v8_1[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[11] simplest_analog_switch_ena1v8_1[1]/avdd simplest_analog_switch_ena1v8_1[1]/dvdd
+ simplest_analog_switch_ena1v8_1[1]/avss simplest_analog_switch_ena1v8_0[11]/on simplest_analog_switch_ena1v8_1[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[12] simplest_analog_switch_ena1v8_1[2]/avdd simplest_analog_switch_ena1v8_1[2]/dvdd
+ simplest_analog_switch_ena1v8_1[2]/avss simplest_analog_switch_ena1v8_0[12]/on simplest_analog_switch_ena1v8_1[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[2]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[13] simplest_analog_switch_ena1v8_1[3]/avdd simplest_analog_switch_ena1v8_1[3]/dvdd
+ simplest_analog_switch_ena1v8_1[3]/avss simplest_analog_switch_ena1v8_0[13]/on simplest_analog_switch_ena1v8_1[3]/out
+ VSUBS simplest_analog_switch_ena1v8_6[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[14] simplest_analog_switch_ena1v8_0[14]/avdd simplest_analog_switch_ena1v8_0[14]/dvdd
+ simplest_analog_switch_ena1v8_0[14]/avss simplest_analog_switch_ena1v8_0[14]/on
+ simplest_analog_switch_ena1v8_1[3]/out VSUBS simplest_analog_switch_ena1v8_6[1]/in
+ simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[15] simplest_analog_switch_ena1v8_5[0]/avdd simplest_analog_switch_ena1v8_5[0]/dvdd
+ simplest_analog_switch_ena1v8_5[0]/avss simplest_analog_switch_ena1v8_0[15]/on simplest_analog_switch_ena1v8_5[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[5]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[16] simplest_analog_switch_ena1v8_5[1]/avdd simplest_analog_switch_ena1v8_5[1]/dvdd
+ simplest_analog_switch_ena1v8_5[1]/avss simplest_analog_switch_ena1v8_0[16]/on simplest_analog_switch_ena1v8_5[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[6]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[17] simplest_analog_switch_ena1v8_5[2]/avdd simplest_analog_switch_ena1v8_5[2]/dvdd
+ simplest_analog_switch_ena1v8_5[2]/avss simplest_analog_switch_ena1v8_0[17]/on simplest_analog_switch_ena1v8_5[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[7]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[18] simplest_analog_switch_ena1v8_5[3]/avdd simplest_analog_switch_ena1v8_5[3]/dvdd
+ simplest_analog_switch_ena1v8_5[3]/avss simplest_analog_switch_ena1v8_0[18]/on simplest_analog_switch_ena1v8_5[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[8]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[19] simplest_analog_switch_ena1v8_0[19]/avdd simplest_analog_switch_ena1v8_0[19]/dvdd
+ simplest_analog_switch_ena1v8_0[19]/avss simplest_analog_switch_ena1v8_0[19]/on
+ simplest_analog_switch_ena1v8_5[3]/out VSUBS simplest_analog_switch_ena1v8_4[0]/in
+ simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[20] simplest_analog_switch_ena1v8_6[0]/avdd simplest_analog_switch_ena1v8_6[0]/dvdd
+ simplest_analog_switch_ena1v8_6[0]/avss simplest_analog_switch_ena1v8_0[20]/on simplest_analog_switch_ena1v8_6[2]/out
+ VSUBS simplest_analog_switch_ena1v8_0[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[21] simplest_analog_switch_ena1v8_6[1]/avdd simplest_analog_switch_ena1v8_6[1]/dvdd
+ simplest_analog_switch_ena1v8_6[1]/avss simplest_analog_switch_ena1v8_0[21]/on simplest_analog_switch_ena1v8_6[2]/out
+ VSUBS simplest_analog_switch_ena1v8_0[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[22] simplest_analog_switch_ena1v8_6[2]/avdd simplest_analog_switch_ena1v8_6[2]/dvdd
+ simplest_analog_switch_ena1v8_6[2]/avss simplest_analog_switch_ena1v8_0[22]/on simplest_analog_switch_ena1v8_6[2]/out
+ VSUBS simplest_analog_switch_ena1v8_0[2]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[23] simplest_analog_switch_ena1v8_0[23]/avdd simplest_analog_switch_ena1v8_0[23]/dvdd
+ simplest_analog_switch_ena1v8_0[23]/avss simplest_analog_switch_ena1v8_0[23]/on
+ simplest_analog_switch_ena1v8_6[2]/out VSUBS simplest_analog_switch_ena1v8_2[0]/in
+ simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[24] simplest_analog_switch_ena1v8_7[0]/avdd simplest_analog_switch_ena1v8_7[0]/dvdd
+ simplest_analog_switch_ena1v8_7[0]/avss simplest_analog_switch_ena1v8_0[24]/on simplest_analog_switch_ena1v8_7[1]/out
+ VSUBS simplest_analog_switch_ena1v8_0[5]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[25] simplest_analog_switch_ena1v8_7[1]/avdd simplest_analog_switch_ena1v8_7[1]/dvdd
+ simplest_analog_switch_ena1v8_7[1]/avss simplest_analog_switch_ena1v8_0[25]/on simplest_analog_switch_ena1v8_7[1]/out
+ VSUBS simplest_analog_switch_ena1v8_0[6]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[26] simplest_analog_switch_ena1v8_0[26]/avdd simplest_analog_switch_ena1v8_0[26]/dvdd
+ simplest_analog_switch_ena1v8_0[26]/avss simplest_analog_switch_ena1v8_0[26]/on
+ simplest_analog_switch_ena1v8_7[1]/out VSUBS simplest_analog_switch_ena1v8_0[7]/in
+ simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[27] simplest_analog_switch_ena1v8_4[0]/avdd simplest_analog_switch_ena1v8_4[0]/dvdd
+ simplest_analog_switch_ena1v8_4[0]/avss simplest_analog_switch_ena1v8_0[27]/on simplest_analog_switch_ena1v8_4[1]/out
+ VSUBS simplest_analog_switch_ena1v8_0[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[28] simplest_analog_switch_ena1v8_4[1]/avdd simplest_analog_switch_ena1v8_4[1]/dvdd
+ simplest_analog_switch_ena1v8_4[1]/avss simplest_analog_switch_ena1v8_0[28]/on simplest_analog_switch_ena1v8_4[1]/out
+ VSUBS simplest_analog_switch_ena1v8_0[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[29] simplest_analog_switch_ena1v8_0[29]/avdd simplest_analog_switch_ena1v8_0[29]/dvdd
+ simplest_analog_switch_ena1v8_0[29]/avss simplest_analog_switch_ena1v8_0[29]/on
+ simplest_analog_switch_ena1v8_4[1]/out VSUBS simplest_analog_switch_ena1v8_0[2]/in
+ simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[0] simplest_analog_switch_ena1v8_1[0]/avdd simplest_analog_switch_ena1v8_1[0]/dvdd
+ simplest_analog_switch_ena1v8_1[0]/avss simplest_analog_switch_ena1v8_1[0]/on simplest_analog_switch_ena1v8_1[3]/out
+ VSUBS simplest_analog_switch_ena1v8_2[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1] simplest_analog_switch_ena1v8_1[1]/avdd simplest_analog_switch_ena1v8_1[1]/dvdd
+ simplest_analog_switch_ena1v8_1[1]/avss simplest_analog_switch_ena1v8_1[1]/on simplest_analog_switch_ena1v8_1[3]/out
+ VSUBS simplest_analog_switch_ena1v8_2[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[2] simplest_analog_switch_ena1v8_1[2]/avdd simplest_analog_switch_ena1v8_1[2]/dvdd
+ simplest_analog_switch_ena1v8_1[2]/avss simplest_analog_switch_ena1v8_1[2]/on simplest_analog_switch_ena1v8_1[3]/out
+ VSUBS simplest_analog_switch_ena1v8_6[2]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[3] simplest_analog_switch_ena1v8_1[3]/avdd simplest_analog_switch_ena1v8_1[3]/dvdd
+ simplest_analog_switch_ena1v8_1[3]/avss simplest_analog_switch_ena1v8_1[3]/on simplest_analog_switch_ena1v8_1[3]/out
+ VSUBS simplest_analog_switch_ena1v8_2[3]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_2[0] simplest_analog_switch_ena1v8_2[0]/avdd simplest_analog_switch_ena1v8_2[0]/dvdd
+ simplest_analog_switch_ena1v8_2[0]/avss simplest_analog_switch_ena1v8_2[0]/on simplest_analog_switch_ena1v8_2[3]/out
+ VSUBS simplest_analog_switch_ena1v8_2[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_2[1] simplest_analog_switch_ena1v8_2[1]/avdd simplest_analog_switch_ena1v8_2[1]/dvdd
+ simplest_analog_switch_ena1v8_2[1]/avss simplest_analog_switch_ena1v8_2[1]/on simplest_analog_switch_ena1v8_2[3]/out
+ VSUBS simplest_analog_switch_ena1v8_2[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_2[2] simplest_analog_switch_ena1v8_2[2]/avdd simplest_analog_switch_ena1v8_2[2]/dvdd
+ simplest_analog_switch_ena1v8_2[2]/avss simplest_analog_switch_ena1v8_2[2]/on simplest_analog_switch_ena1v8_2[3]/out
+ VSUBS simplest_analog_switch_ena1v8_6[2]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_2[3] simplest_analog_switch_ena1v8_2[3]/avdd simplest_analog_switch_ena1v8_2[3]/dvdd
+ simplest_analog_switch_ena1v8_2[3]/avss simplest_analog_switch_ena1v8_2[3]/on simplest_analog_switch_ena1v8_2[3]/out
+ VSUBS simplest_analog_switch_ena1v8_2[3]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_3[0] simplest_analog_switch_ena1v8_3[0]/avdd simplest_analog_switch_ena1v8_3[0]/dvdd
+ simplest_analog_switch_ena1v8_3[0]/avss simplest_analog_switch_ena1v8_3[0]/on simplest_analog_switch_ena1v8_3[3]/out
+ VSUBS simplest_analog_switch_ena1v8_5[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_3[1] simplest_analog_switch_ena1v8_3[1]/avdd simplest_analog_switch_ena1v8_3[1]/dvdd
+ simplest_analog_switch_ena1v8_3[1]/avss simplest_analog_switch_ena1v8_3[1]/on simplest_analog_switch_ena1v8_3[3]/out
+ VSUBS simplest_analog_switch_ena1v8_7[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_3[2] simplest_analog_switch_ena1v8_3[2]/avdd simplest_analog_switch_ena1v8_3[2]/dvdd
+ simplest_analog_switch_ena1v8_3[2]/avss simplest_analog_switch_ena1v8_3[2]/on simplest_analog_switch_ena1v8_3[3]/out
+ VSUBS simplest_analog_switch_ena1v8_5[2]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_3[3] simplest_analog_switch_ena1v8_3[3]/avdd simplest_analog_switch_ena1v8_3[3]/dvdd
+ simplest_analog_switch_ena1v8_3[3]/avss simplest_analog_switch_ena1v8_3[3]/on simplest_analog_switch_ena1v8_3[3]/out
+ VSUBS simplest_analog_switch_ena1v8_7[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_4[0] simplest_analog_switch_ena1v8_4[0]/avdd simplest_analog_switch_ena1v8_4[0]/dvdd
+ simplest_analog_switch_ena1v8_4[0]/avss simplest_analog_switch_ena1v8_4[0]/on simplest_analog_switch_ena1v8_4[1]/out
+ VSUBS simplest_analog_switch_ena1v8_4[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_4[1] simplest_analog_switch_ena1v8_4[1]/avdd simplest_analog_switch_ena1v8_4[1]/dvdd
+ simplest_analog_switch_ena1v8_4[1]/avss simplest_analog_switch_ena1v8_4[1]/on simplest_analog_switch_ena1v8_4[1]/out
+ VSUBS simplest_analog_switch_ena1v8_5[2]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_5[0] simplest_analog_switch_ena1v8_5[0]/avdd simplest_analog_switch_ena1v8_5[0]/dvdd
+ simplest_analog_switch_ena1v8_5[0]/avss simplest_analog_switch_ena1v8_5[0]/on simplest_analog_switch_ena1v8_5[3]/out
+ VSUBS simplest_analog_switch_ena1v8_5[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_5[1] simplest_analog_switch_ena1v8_5[1]/avdd simplest_analog_switch_ena1v8_5[1]/dvdd
+ simplest_analog_switch_ena1v8_5[1]/avss simplest_analog_switch_ena1v8_5[1]/on simplest_analog_switch_ena1v8_5[3]/out
+ VSUBS simplest_analog_switch_ena1v8_7[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_5[2] simplest_analog_switch_ena1v8_5[2]/avdd simplest_analog_switch_ena1v8_5[2]/dvdd
+ simplest_analog_switch_ena1v8_5[2]/avss simplest_analog_switch_ena1v8_5[2]/on simplest_analog_switch_ena1v8_5[3]/out
+ VSUBS simplest_analog_switch_ena1v8_5[2]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_5[3] simplest_analog_switch_ena1v8_5[3]/avdd simplest_analog_switch_ena1v8_5[3]/dvdd
+ simplest_analog_switch_ena1v8_5[3]/avss simplest_analog_switch_ena1v8_5[3]/on simplest_analog_switch_ena1v8_5[3]/out
+ VSUBS simplest_analog_switch_ena1v8_7[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_6[0] simplest_analog_switch_ena1v8_6[0]/avdd simplest_analog_switch_ena1v8_6[0]/dvdd
+ simplest_analog_switch_ena1v8_6[0]/avss simplest_analog_switch_ena1v8_6[0]/on simplest_analog_switch_ena1v8_6[2]/out
+ VSUBS simplest_analog_switch_ena1v8_6[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_6[1] simplest_analog_switch_ena1v8_6[1]/avdd simplest_analog_switch_ena1v8_6[1]/dvdd
+ simplest_analog_switch_ena1v8_6[1]/avss simplest_analog_switch_ena1v8_6[1]/on simplest_analog_switch_ena1v8_6[2]/out
+ VSUBS simplest_analog_switch_ena1v8_6[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_6[2] simplest_analog_switch_ena1v8_6[2]/avdd simplest_analog_switch_ena1v8_6[2]/dvdd
+ simplest_analog_switch_ena1v8_6[2]/avss simplest_analog_switch_ena1v8_6[2]/on simplest_analog_switch_ena1v8_6[2]/out
+ VSUBS simplest_analog_switch_ena1v8_6[2]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_7[0] simplest_analog_switch_ena1v8_7[0]/avdd simplest_analog_switch_ena1v8_7[0]/dvdd
+ simplest_analog_switch_ena1v8_7[0]/avss simplest_analog_switch_ena1v8_7[0]/on simplest_analog_switch_ena1v8_7[1]/out
+ VSUBS simplest_analog_switch_ena1v8_7[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_7[1] simplest_analog_switch_ena1v8_7[1]/avdd simplest_analog_switch_ena1v8_7[1]/dvdd
+ simplest_analog_switch_ena1v8_7[1]/avss simplest_analog_switch_ena1v8_7[1]/on simplest_analog_switch_ena1v8_7[1]/out
+ VSUBS simplest_analog_switch_ena1v8_7[1]/in simplest_analog_switch_ena1v8
.ends

.subckt simple_switch_array_16 vdda0 simplest_analog_switch_ena1v8_1[1|1]/on left_lp_opamp_p
+ comp_p simplest_analog_switch_ena1v8_1[3|3]/on left_lp_opamp_n simplest_analog_switch_ena1v8_1[0|1]/on
+ comp_n simplest_analog_switch_ena1v8_1[1|0]/on simplest_analog_switch_ena1v8_1[2|1]/on
+ simplest_analog_switch_ena1v8_1[3|2]/on simplest_analog_switch_ena1v8_1[0|2]/on
+ simplest_analog_switch_ena1v8_1[1|3]/on right_hgbw_opamp_p simplest_analog_switch_ena1v8_1[0|3]/on
+ right_hgbw_opamp_n left_hgbw_opamp_p left_hgbw_opamp_n simplest_analog_switch_ena1v8_1[2|3]/on
+ simplest_analog_switch_ena1v8_1[2|0]/on right_instramp_p simplest_analog_switch_ena1v8_1[3|1]/on
+ right_instramp_n ulpcomp_p simplest_analog_switch_ena1v8_1[2|2]/on ulpcomp_n sio1
+ right_lp_opamp_p sio0 simplest_analog_switch_ena1v8_1[1|2]/on left_instramp_p right_lp_opamp_n
+ vccd0 simplest_analog_switch_ena1v8_1[3|0]/on left_instramp_n simplest_analog_switch_ena1v8_1[0|0]/on
+ vssa0 vssd0
Xsimplest_analog_switch_ena1v8_1[0|0] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[0|0]/on
+ sio1 vssd0 ulpcomp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1|0] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[1|0]/on
+ sio1 vssd0 comp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[2|0] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[2|0]/on
+ sio0 vssd0 ulpcomp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[3|0] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[3|0]/on
+ sio0 vssd0 comp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[0|1] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[0|1]/on
+ sio1 vssd0 left_lp_opamp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1|1] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[1|1]/on
+ sio1 vssd0 left_instramp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[2|1] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[2|1]/on
+ sio0 vssd0 left_lp_opamp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[3|1] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[3|1]/on
+ sio0 vssd0 left_instramp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[0|2] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[0|2]/on
+ sio1 vssd0 right_hgbw_opamp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1|2] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[1|2]/on
+ sio1 vssd0 left_hgbw_opamp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[2|2] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[2|2]/on
+ sio0 vssd0 right_hgbw_opamp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[3|2] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[3|2]/on
+ sio0 vssd0 left_hgbw_opamp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[0|3] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[0|3]/on
+ sio1 vssd0 right_instramp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1|3] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[1|3]/on
+ sio1 vssd0 right_lp_opamp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[2|3] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[2|3]/on
+ sio0 vssd0 right_instramp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[3|3] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[3|3]/on
+ sio0 vssd0 right_lp_opamp_p simplest_analog_switch_ena1v8
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_KB5CJD m4_n1349_n1080# c2_n1269_n1000#
X0 c2_n1269_n1000# m4_n1349_n1080# sky130_fd_pr__cap_mim_m3_2 l=10 w=10
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_C3WBNQ a_n296_n522# a_n158_n300# a_n100_n388#
+ a_100_n300#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n296_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RK a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_QRKT8P a_n296_n522# a_n158_n300# a_n100_n388#
+ a_100_n300#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n296_n522# sky130_fd_pr__nfet_05v0_nvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ZMKT8P a_n296_n522# a_n158_n300# a_n100_n388#
+ a_100_n300#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n296_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt bias_nstack itail ena nbias avss vcasc
XXM12 avss avss nbias m1_3726_n2502# sky130_fd_pr__nfet_g5v0d10v5_C3WBNQ
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RK_0 avss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RK
XXM6 avss vcasc nbias m1_3726_n2502# sky130_fd_pr__nfet_05v0_nvt_QRKT8P
XXM7 avss vcasc ena itail sky130_fd_pr__nfet_g5v0d10v5_ZMKT8P
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RJ a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__res_high_po_0p35_P35QVK a_380_2984# a_5692_n3416# a_n3770_2984#
+ a_3866_2984# a_3202_n3416# a_n1446_n3416# a_n284_n3416# a_n616_2984# a_4696_n3416#
+ a_4198_2984# a_2206_n3416# a_n1114_2984# a_n4102_2984# a_n616_n3416# a_6190_n3416#
+ a_n6592_2984# a_2372_2984# a_n5762_n3416# a_5360_2984# a_214_2984# a_n3604_2984#
+ a_1210_n3416# a_5194_n3416# a_6522_n3416# a_n4766_n3416# a_1874_2984# a_4862_2984#
+ a_4198_n3416# a_5526_n3416# a_5194_2984# a_n6260_n3416# a_878_n3416# a_n3438_2984#
+ a_n2110_2984# a_n6426_2984# a_2206_2984# a_n118_n3416# a_n3770_n3416# a_4696_2984#
+ a_n5264_n3416# a_48_2984# a_4530_n3416# a_n2774_n3416# a_n1612_2984# a_n4600_2984#
+ a_n5928_2984# a_1708_2984# a_6024_n3416# a_n4268_n3416# a_2870_2984# a_3534_n3416#
+ a_712_2984# a_n1778_n3416# a_5028_2984# a_5028_n3416# a_n948_2984# a_2538_n3416#
+ a_6190_2984# a_n1446_2984# a_n3272_n3416# a_n4434_2984# a_n4600_n3416# a_3202_2984#
+ a_n948_n3416# a_5692_2984# a_380_n3416# a_546_2984# a_4032_n3416# a_n2276_n3416#
+ a_n3604_n3416# a_n3936_2984# a_1542_n3416# a_2704_2984# a_3036_n3416# a_712_n3416#
+ a_n2608_n3416# a_n4268_2984# a_3036_2984# a_6024_2984# a_5858_n3416# a_n1280_n3416#
+ a_n6592_n3416# a_n2442_2984# a_n4102_n3416# a_2538_2984# a_n5430_2984# a_2040_n3416#
+ a_5526_2984# a_1210_2984# a_n1612_n3416# a_n5596_n3416# a_4862_n3416# a_n450_n3416#
+ a_n1944_2984# a_n3106_n3416# a_n4932_2984# a_1044_n3416# a_n450_2984# a_3700_2984#
+ a_6356_n3416# a_214_n3416# a_n5928_n3416# a_n6722_n3546# a_3866_n3416# a_n2276_2984#
+ a_n5264_2984# a_1044_2984# a_4032_2984# a_n2110_n3416# a_n6094_n3416# a_n1778_2984#
+ a_n4766_2984# a_5360_n3416# a_n284_2984# a_3534_2984# a_n4932_n3416# a_6522_2984#
+ a_n1114_n3416# a_2870_n3416# a_n5098_n3416# a_n6426_n3416# a_878_2984# a_4364_n3416#
+ a_n5098_2984# a_n3936_n3416# a_n2940_2984# a_1874_n3416# a_3368_n3416# a_n3272_2984#
+ a_3368_2984# a_48_n3416# a_n6260_2984# a_2040_2984# a_6356_2984# a_n5430_n3416#
+ a_n2940_n3416# a_n118_2984# a_n2774_2984# a_n4434_n3416# a_n5762_2984# a_1542_2984#
+ a_2372_n3416# a_4530_2984# a_5858_2984# a_3700_n3416# a_n1944_n3416# a_n3438_n3416#
+ a_n6094_2984# a_n782_n3416# a_1376_n3416# a_n782_2984# a_2704_n3416# a_546_n3416#
+ a_n3106_2984# a_n1280_2984# a_n5596_2984# a_1376_2984# a_1708_n3416# a_4364_2984#
+ a_n2442_n3416# a_n2608_2984#
X0 a_n3936_2984# a_n3936_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X1 a_n1612_2984# a_n1612_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X2 a_n450_2984# a_n450_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X3 a_n284_2984# a_n284_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X4 a_n4434_2984# a_n4434_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X5 a_48_2984# a_48_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X6 a_n6592_2984# a_n6592_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X7 a_2704_2984# a_2704_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X8 a_4862_2984# a_4862_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X9 a_3202_2984# a_3202_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X10 a_5360_2984# a_5360_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X11 a_5526_2984# a_5526_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X12 a_n948_2984# a_n948_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X13 a_n782_2984# a_n782_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X14 a_6024_2984# a_6024_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X15 a_n4932_2984# a_n4932_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X16 a_1376_2984# a_1376_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X17 a_878_2984# a_878_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X18 a_4198_2984# a_4198_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X19 a_3700_2984# a_3700_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X20 a_n3770_2984# a_n3770_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X21 a_n1446_2984# a_n1446_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X22 a_6522_2984# a_6522_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X23 a_n4268_2984# a_n4268_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X24 a_n2110_2984# a_n2110_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X25 a_1874_2984# a_1874_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X26 a_2372_2984# a_2372_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X27 a_2538_2984# a_2538_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X28 a_4696_2984# a_4696_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X29 a_3036_2984# a_3036_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X30 a_5194_2984# a_5194_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X31 a_n1944_2984# a_n1944_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X32 a_n4766_2984# a_n4766_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X33 a_n2608_2984# a_n2608_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X34 a_n2442_2984# a_n2442_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X35 a_214_2984# a_214_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X36 a_n5430_2984# a_n5430_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X37 a_n5264_2984# a_n5264_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X38 a_n3106_2984# a_n3106_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X39 a_2870_2984# a_2870_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X40 a_n1280_2984# a_n1280_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X41 a_1210_2984# a_1210_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X42 a_3534_2984# a_3534_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X43 a_5692_2984# a_5692_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X44 a_5858_2984# a_5858_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X45 a_712_2984# a_712_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X46 a_4032_2984# a_4032_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X47 a_6190_2984# a_6190_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X48 a_6356_2984# a_6356_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X49 a_n118_2984# a_n118_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X50 a_n5928_2984# a_n5928_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X51 a_n5762_2984# a_n5762_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X52 a_n3604_2984# a_n3604_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X53 a_n6426_2984# a_n6426_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X54 a_n4102_2984# a_n4102_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X55 a_n1778_2984# a_n1778_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X56 a_n4600_2984# a_n4600_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X57 a_n2276_2984# a_n2276_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X58 a_4530_2984# a_4530_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X59 a_n5098_2984# a_n5098_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X60 a_n616_2984# a_n616_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X61 a_1044_2984# a_1044_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X62 a_3368_2984# a_3368_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X63 a_380_2984# a_380_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X64 a_546_2984# a_546_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X65 a_n2940_2984# a_n2940_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X66 a_n2774_2984# a_n2774_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X67 a_n5596_2984# a_n5596_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X68 a_n3438_2984# a_n3438_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X69 a_n3272_2984# a_n3272_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X70 a_n1114_2984# a_n1114_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X71 a_n6260_2984# a_n6260_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X72 a_n6094_2984# a_n6094_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X73 a_1542_2984# a_1542_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X74 a_1708_2984# a_1708_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X75 a_3866_2984# a_3866_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X76 a_2040_2984# a_2040_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X77 a_2206_2984# a_2206_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X78 a_4364_2984# a_4364_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X79 a_5028_2984# a_5028_n3416# a_n6722_n3546# sky130_fd_pr__res_high_po_0p35 l=30
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ a_n158_n300# w_n362_n597# a_n100_n397#
+ a_100_n300#
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n362_n597# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_H75TTW a_n158_n300# w_n362_n597# a_n100_n397#
+ a_100_n300#
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n362_n597# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt bias_pstack pcasc enb itail vcasc pbias avss avdd
XXM13 m1_2150_n1558# avdd pcasc vcasc sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ
Xsky130_fd_pr__pfet_g5v0d10v5_G8LMTZ_0 itail avdd enb vcasc sky130_fd_pr__pfet_g5v0d10v5_G8LMTZ
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RK_0 avss enb sky130_fd_pr__diode_pw2nd_05v5_FT76RK
Xsky130_fd_pr__pfet_g5v0d10v5_H75TTW_0 m1_2150_n1558# avdd pbias avdd sky130_fd_pr__pfet_g5v0d10v5_H75TTW
.ends

.subckt sky130_fd_pr__res_high_po_0p35_L4QTBM a_3451_2984# a_4447_n3416# a_795_2984#
+ a_1957_n3416# a_n5181_n3416# a_n201_2984# a_n2691_n3416# a_2953_2984# a_n2027_2984#
+ a_n4185_n3416# a_n5015_2984# a_n5513_n3416# a_3451_n3416# a_n1695_n3416# a_3285_2984#
+ a_n3189_n3416# a_n1529_2984# a_n4517_n3416# a_n4517_2984# a_2455_n3416# a_297_n3416#
+ a_n2691_2984# a_2787_2984# a_629_2984# a_n35_2984# a_n865_n3416# a_1459_n3416# a_629_n3416#
+ a_n2193_n3416# a_n3521_n3416# a_n3023_2984# a_n5015_n3416# a_3119_2984# a_n1197_n3416#
+ a_n2525_n3416# a_1293_2984# a_4281_2984# a_n4019_n3416# a_n2525_2984# a_n5513_2984#
+ a_n1529_n3416# a_3783_2984# a_4779_n3416# a_n367_n3416# a_n533_2984# a_n3023_n3416#
+ a_n2359_2984# a_131_n3416# a_n1031_2984# a_n5347_2984# a_1127_2984# a_4115_2984#
+ a_n2027_n3416# a_3783_n3416# a_5277_n3416# a_131_2984# a_n4849_n3416# a_n4849_2984#
+ a_n367_2984# a_n3521_2984# a_n5643_n3546# a_2787_n3416# a_3617_2984# a_1791_2984#
+ a_n1031_n3416# a_4281_n3416# a_n3853_n3416# a_1791_n3416# a_n3355_2984# a_n5347_n3416#
+ a_961_n3416# a_2123_2984# a_3285_n3416# a_4613_n3416# a_5111_2984# a_n201_n3416#
+ a_n2857_n3416# a_n2857_2984# a_2289_n3416# a_1625_2984# a_3617_n3416# a_4613_2984#
+ a_n4351_n3416# a_n699_n3416# a_n3189_2984# a_n1861_n3416# a_n865_2984# a_5111_n3416#
+ a_n3355_n3416# a_1293_n3416# a_2621_n3416# a_n1363_2984# a_n4351_2984# a_463_n3416#
+ a_1459_2984# a_4115_n3416# a_4447_2984# a_n2359_n3416# a_463_2984# a_1625_n3416#
+ a_n699_2984# a_n3853_2984# a_3119_n3416# a_3949_2984# a_2621_2984# a_n1197_2984#
+ a_n1363_n3416# a_n4185_2984# a_297_2984# a_2123_n3416# a_n3687_2984# a_2455_2984#
+ a_5443_2984# a_n533_n3416# a_4945_n3416# a_1127_n3416# a_n1861_2984# a_1957_2984#
+ a_3949_n3416# a_4945_2984# a_n35_n3416# a_n4019_2984# a_n4683_n3416# a_961_2984#
+ a_n2193_2984# a_2289_2984# a_n5181_2984# a_5277_2984# a_5443_n3416# a_n3687_n3416#
+ a_2953_n3416# a_n1695_2984# a_n4683_2984# a_795_n3416# a_4779_2984#
X0 a_2953_2984# a_2953_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X1 a_n1197_2984# a_n1197_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X2 a_3451_2984# a_3451_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X3 a_3617_2984# a_3617_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X4 a_4115_2984# a_4115_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X5 a_2289_2984# a_2289_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X6 a_n3521_2984# a_n3521_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X7 a_n2359_2984# a_n2359_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X8 a_n1695_2984# a_n1695_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X9 a_4613_2984# a_4613_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X10 a_n2193_2984# a_n2193_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X11 a_5111_2984# a_5111_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X12 a_n533_2984# a_n533_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X13 a_2787_2984# a_2787_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X14 a_1127_2984# a_1127_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X15 a_3285_2984# a_3285_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X16 a_463_2984# a_463_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X17 a_629_2984# a_629_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X18 a_n2857_2984# a_n2857_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X19 a_n2691_2984# a_n2691_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X20 a_n3355_2984# a_n3355_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X21 a_n1031_2984# a_n1031_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X22 a_n4019_2984# a_n4019_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X23 a_n35_2984# a_n35_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X24 a_1625_2984# a_1625_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X25 a_3949_2984# a_3949_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X26 a_2123_2984# a_2123_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X27 a_3783_2984# a_3783_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X28 a_4447_2984# a_4447_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X29 a_961_2984# a_961_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X30 a_4281_2984# a_4281_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X31 a_n367_2984# a_n367_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X32 a_n4517_2984# a_n4517_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X33 a_n3853_2984# a_n3853_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X34 a_n5015_2984# a_n5015_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X35 a_n4351_2984# a_n4351_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X36 a_297_2984# a_297_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X37 a_2621_2984# a_2621_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X38 a_4945_2984# a_4945_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X39 a_n3189_2984# a_n3189_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X40 a_5443_2984# a_5443_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X41 a_n865_2984# a_n865_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X42 a_1293_2984# a_1293_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X43 a_1459_2984# a_1459_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X44 a_n5513_2984# a_n5513_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X45 a_795_2984# a_795_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X46 a_n3687_2984# a_n3687_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X47 a_n1529_2984# a_n1529_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X48 a_n1363_2984# a_n1363_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X49 a_n4185_2984# a_n4185_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X50 a_n2027_2984# a_n2027_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X51 a_1791_2984# a_1791_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X52 a_1957_2984# a_1957_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X53 a_n201_2984# a_n201_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X54 a_2455_2984# a_2455_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X55 a_4779_2984# a_4779_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X56 a_3119_2984# a_3119_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X57 a_5277_2984# a_5277_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X58 a_n1861_2984# a_n1861_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X59 a_n699_2984# a_n699_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X60 a_n4849_2984# a_n4849_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X61 a_n4683_2984# a_n4683_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X62 a_n2525_2984# a_n2525_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X63 a_131_2984# a_131_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X64 a_n5347_2984# a_n5347_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X65 a_n5181_2984# a_n5181_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
X66 a_n3023_2984# a_n3023_n3416# a_n5643_n3546# sky130_fd_pr__res_high_po_0p35 l=30
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_F3TL5C a_100_n200# a_n292_n422# a_n158_n200# a_n100_n288#
X0 a_100_n200# a_n100_n288# a_n158_n200# a_n292_n422# sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_56WC32 a_100_n200# a_n158_n200# a_n332_n422#
+ a_n100_n288#
X0 a_100_n200# a_n100_n288# a_n158_n200# a_n332_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QSDYAY w_n487_n497# a_29_n297# a_n287_n200# a_n229_n297#
+ a_229_n200# a_n29_n200#
X0 a_n29_n200# a_n229_n297# a_n287_n200# w_n487_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X1 a_229_n200# a_29_n297# a_n29_n200# w_n487_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_V5WCXY a_n287_n200# a_n487_n288# a_229_n200#
+ a_n545_n200# a_29_n288# a_487_n200# a_n29_n200# a_n229_n288# a_287_n288# a_n679_n422#
X0 a_n29_n200# a_n229_n288# a_n287_n200# a_n679_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_229_n200# a_29_n288# a_n29_n200# a_n679_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_n287_n200# a_n487_n288# a_n545_n200# a_n679_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X3 a_487_n200# a_287_n288# a_229_n200# a_n679_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt bias_amp nbias ena inp inn out avss avdd
Xsky130_fd_pr__nfet_05v0_nvt_F3TL5C_0 m1_5615_3673# avss m1_7291_3557# ena sky130_fd_pr__nfet_05v0_nvt_F3TL5C
Xsky130_fd_pr__nfet_g5v0d10v5_56WC32_0 m1_7291_3557# avss avss nbias sky130_fd_pr__nfet_g5v0d10v5_56WC32
Xsky130_fd_pr__pfet_g5v0d10v5_QSDYAY_0 avdd m1_6016_4428# m1_6016_4428# m1_6016_4428#
+ out avdd sky130_fd_pr__pfet_g5v0d10v5_QSDYAY
Xsky130_fd_pr__nfet_g5v0d10v5_V5WCXY_0 m1_6016_4428# inp out m1_5615_3673# inn m1_5615_3673#
+ m1_5615_3673# inp inn avss sky130_fd_pr__nfet_g5v0d10v5_V5WCXY
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MQZGVK m3_n686_n2520# c1_n646_n2480#
X0 c1_n646_n2480# m3_n686_n2520# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
X1 c1_n646_n2480# m3_n686_n2520# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
X2 c1_n646_n2480# m3_n686_n2520# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
X3 c1_n646_n2480# m3_n686_n2520# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
.ends

.subckt bias_generator_fe snk_test0 src_test0 vbg ref_in ena_snk_test0 ena_src_test0
+ ref_sel_vbg dvdd dvss bias_amp_0/out avdd bias_amp_0/nbias ena bias_pstack_0[9]/pcasc
+ avss
Xbias_nstack_0[0] snk_test0 ena_test0_3v3 bias_amp_0/nbias avss bias_nstack_0[0]/vcasc
+ bias_nstack
Xbias_nstack_0[1] snk_test0 ena_test0_3v3 bias_amp_0/nbias avss bias_nstack_0[1]/vcasc
+ bias_nstack
Xbias_nstack_0[2] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[3] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[4] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[5] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[6] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[7] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[8] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[9] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[10] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[11] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[12] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[13] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[14] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[15] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[16] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[17] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[18] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[19] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[20] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[21] bias_nstack_0[9]/itail ena_3v3 bias_amp_0/nbias avss bias_amp_0/nbias
+ bias_nstack
Xbias_nstack_0[22] bias_amp_0/out enb_vbg_3v3 bias_amp_0/nbias avss bias_nstack_0[22]/vcasc
+ bias_nstack
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0 avss vbg sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
XXR2 m1_26761_7166# m1_31907_766# m1_22445_7166# m1_30081_7166# m1_29583_766# m1_24935_766#
+ m1_25931_766# m1_25765_7166# m1_30911_766# m1_30413_7166# m1_28587_766# m1_25101_7166#
+ m1_22113_7166# m1_25599_766# m1_32571_766# m1_19789_7166# m1_28753_7166# m1_20619_766#
+ m1_31741_7166# m1_26429_7166# m1_22777_7166# m1_27591_766# m1_31575_766# bias_nstack_0[9]/itail
+ m1_21615_766# m1_28089_7166# m1_31077_7166# m1_30579_766# m1_31907_766# m1_31409_7166#
+ m1_19955_766# m1_27259_766# m1_22777_7166# m1_24105_7166# m1_19789_7166# m1_28421_7166#
+ m1_26263_766# m1_22611_766# m1_31077_7166# m1_20951_766# m1_26429_7166# m1_30911_766#
+ m1_23607_766# m1_24769_7166# m1_21781_7166# m1_20453_7166# m1_28089_7166# m1_32239_766#
+ m1_21947_766# m1_29085_7166# m1_29915_766# m1_27093_7166# m1_24603_766# m1_31409_7166#
+ m1_31243_766# m1_25433_7166# m1_28919_766# m1_32405_7166# m1_24769_7166# m1_22943_766#
+ m1_21781_7166# m1_21615_766# m1_29417_7166# m1_25267_766# m1_32073_7166# m1_26595_766#
+ m1_26761_7166# m1_30247_766# m1_23939_766# m1_22611_766# m1_22445_7166# bias_pstack_0[9]/pcasc
+ m1_29085_7166# m1_29251_766# m1_26927_766# m1_23607_766# m1_22113_7166# m1_29417_7166#
+ m1_32405_7166# m1_32239_766# m1_24935_766# ref_in m1_23773_7166# m1_22279_766# m1_28753_7166#
+ m1_20785_7166# m1_28255_766# m1_31741_7166# m1_27425_7166# m1_24603_766# m1_20619_766#
+ m1_31243_766# m1_25931_766# m1_24437_7166# m1_23275_766# m1_21449_7166# m1_27259_766#
+ m1_25765_7166# m1_30081_7166# m1_32571_766# m1_26595_766# m1_20287_766# avss m1_30247_766#
+ m1_24105_7166# m1_21117_7166# m1_27425_7166# m1_30413_7166# m1_24271_766# m1_20287_766#
+ m1_24437_7166# m1_21449_7166# m1_31575_766# m1_26097_7166# m1_29749_7166# m1_21283_766#
+ m1_32737_7166# m1_25267_766# m1_29251_766# m1_21283_766# m1_19955_766# m1_27093_7166#
+ m1_30579_766# m1_21117_7166# m1_22279_766# m1_23441_7166# m1_28255_766# m1_29583_766#
+ m1_23109_7166# m1_29749_7166# m1_26263_766# m1_20121_7166# m1_28421_7166# m1_32737_7166#
+ m1_20951_766# m1_23275_766# m1_26097_7166# m1_23441_7166# m1_21947_766# m1_20453_7166#
+ m1_27757_7166# m1_28587_766# m1_30745_7166# m1_32073_7166# m1_29915_766# m1_24271_766#
+ m1_22943_766# m1_20121_7166# m1_25599_766# m1_27591_766# m1_25433_7166# m1_28919_766#
+ m1_26927_766# m1_23109_7166# m1_25101_7166# m1_20785_7166# m1_27757_7166# bias_pstack_0[9]/pcasc
+ m1_30745_7166# m1_23939_766# m1_23773_7166# sky130_fd_pr__res_high_po_0p35_P35QVK
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0] ena_snk_test0 dvdd dvss avdd avdd ena_test0_3v3
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1] ena_src_test0 dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_2/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[2] ena dvdd dvss avdd avdd ena_3v3 avdd dvss dvss
+ sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[3] ref_sel_vbg dvdd dvss avdd avdd ena_vbg_3v3 avdd
+ dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__inv_2_2 sky130_fd_sc_hvl__inv_2_2/A dvss dvss avdd avdd enb_test0_3v3
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_4 ena_vbg_3v3 dvss dvss avdd avdd enb_vbg_3v3 sky130_fd_sc_hvl__inv_2
Xbias_pstack_0[0] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[0]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[1] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[1]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[2] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[2]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[3] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[3]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[4] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[4]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[5] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[5]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[6] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[6]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[7] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[7]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[8] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[8]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[9] bias_pstack_0[9]/pcasc enb_test0_3v3 src_test0 bias_pstack_0[9]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[10] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[10]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[11] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[11]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[12] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[12]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[13] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[13]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[14] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[14]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[15] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[15]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[16] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[16]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[17] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[17]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[18] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[18]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[19] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[19]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[20] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[20]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[21] bias_pstack_0[9]/pcasc enb_vbg_3v3 bias_amp_0/inp bias_pstack_0[21]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xbias_pstack_0[22] bias_pstack_0[9]/pcasc ena_vbg_3v3 bias_amp_0/out bias_pstack_0[22]/vcasc
+ bias_amp_0/out avss avdd bias_pstack
Xsky130_fd_pr__res_high_po_0p35_L4QTBM_0 m1_17229_7166# m1_18391_766# m1_14573_7166#
+ m1_15735_766# m1_8763_766# m1_13577_7166# m1_11087_766# m1_16897_7166# m1_11917_7166#
+ m1_9759_766# m1_8929_7166# m1_8431_766# m1_17395_766# m1_12083_766# m1_17229_7166#
+ m1_10755_766# m1_12249_7166# m1_9427_766# m1_9261_7166# m1_16399_766# m1_14075_766#
+ m1_11253_7166# m1_16565_7166# m1_14573_7166# m1_13909_7166# m1_13079_766# m1_15403_766#
+ m1_14407_766# m1_11751_766# m1_10423_766# m1_10921_7166# m1_8763_766# m1_16897_7166#
+ m1_12747_766# m1_11419_766# m1_15237_7166# m1_18225_7166# m1_9759_766# m1_11253_7166#
+ bias_amp_0/inp m1_12415_766# m1_17561_7166# m1_18723_766# m1_13411_766# m1_13245_7166#
+ m1_10755_766# m1_11585_7166# m1_14075_766# m1_12913_7166# m1_8597_7166# m1_14905_7166#
+ m1_17893_7166# m1_11751_766# m1_17727_766# m1_19055_766# m1_13909_7166# m1_9095_766#
+ m1_8929_7166# m1_13577_7166# m1_10257_7166# avss m1_16731_766# m1_17561_7166# m1_15569_7166#
+ m1_12747_766# m1_18059_766# m1_10091_766# m1_15735_766# m1_10589_7166# m1_8431_766#
+ m1_14739_766# m1_15901_7166# m1_17063_766# m1_18391_766# m1_18889_7166# m1_13743_766#
+ m1_11087_766# m1_10921_7166# m1_16067_766# m1_15569_7166# m1_17395_766# m1_18557_7166#
+ m1_9427_766# m1_13079_766# m1_10589_7166# m1_12083_766# m1_12913_7166# m1_19055_766#
+ m1_10423_766# m1_15071_766# m1_16399_766# m1_12581_7166# m1_9593_7166# m1_14407_766#
+ m1_15237_7166# m1_18059_766# m1_18225_7166# m1_11419_766# m1_14241_7166# m1_15403_766#
+ m1_13245_7166# m1_9925_7166# m1_17063_766# m1_17893_7166# m1_16565_7166# m1_12581_7166#
+ m1_12415_766# m1_9593_7166# m1_14241_7166# m1_16067_766# m1_10257_7166# m1_16233_7166#
+ m1_19221_7166# m1_13411_766# m1_18723_766# m1_15071_766# m1_11917_7166# m1_15901_7166#
+ m1_17727_766# m1_18889_7166# m1_13743_766# m1_9925_7166# m1_9095_766# m1_14905_7166#
+ m1_11585_7166# m1_16233_7166# m1_8597_7166# m1_19221_7166# avss m1_10091_766# m1_16731_766#
+ m1_12249_7166# m1_9261_7166# m1_14739_766# m1_18557_7166# sky130_fd_pr__res_high_po_0p35_L4QTBM
Xsky130_fd_sc_hvl__diode_2_0 ena dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_11 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_1 ena_snk_test0 dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xbias_amp_0 bias_amp_0/nbias ena_vbg_3v3 bias_amp_0/inp vbg bias_amp_0/out avss avdd
+ bias_amp
Xsky130_fd_sc_hvl__diode_2_2 ena_src_test0 dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_3 ref_sel_vbg dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_pr__cap_mim_m3_1_MQZGVK_0 bias_amp_0/inp bias_amp_0/out sky130_fd_pr__cap_mim_m3_1_MQZGVK
Xsky130_fd_pr__cap_mim_m3_1_MQZGVK_1 bias_amp_0/inp bias_amp_0/out sky130_fd_pr__cap_mim_m3_1_MQZGVK
Xsky130_fd_sc_hvl__decap_4_3 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
.ends

.subckt bias_generator_idac_be avdd dvdd dvss ena[6] ena[3] ena[2] ena[0] ena[1] ena[5]
+ ena[4] ena[7] avss_uq0 avdd_uq0 avdd_uq1 avdd_uq2 a_135144_n10736# m4_89432_13963#
+ a_89514_n1347# m4_89432_n426# a_89514_7744# bias_nstack_3[3]/itail bias_nstack_3[3]/nbias
+ bias_pstack_3[3]/pcasc bias_pstack_2[9]/itail bias_pstack_1[9]/itail bias_pstack_0[9]/itail
+ bias_nstack_1[9]/itail bias_pstack_3[3]/itail avss_uq1 bias_nstack_2[9]/itail bias_nstack_0[9]/itail
+ avss avss_uq2 bias_pstack_3[3]/pbias
Xbias_nstack_0[0] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[0]/vcasc bias_nstack
Xbias_nstack_0[1] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[1]/vcasc bias_nstack
Xbias_nstack_0[2] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[2]/vcasc bias_nstack
Xbias_nstack_0[3] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[3]/vcasc bias_nstack
Xbias_nstack_0[4] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[4]/vcasc bias_nstack
Xbias_nstack_0[5] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[5]/vcasc bias_nstack
Xbias_nstack_0[6] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[6]/vcasc bias_nstack
Xbias_nstack_0[7] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[7]/vcasc bias_nstack
Xbias_nstack_0[8] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[8]/vcasc bias_nstack
Xbias_nstack_0[9] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[9]/vcasc bias_nstack
Xbias_nstack_0[10] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[10]/vcasc bias_nstack
Xbias_nstack_0[11] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[11]/vcasc bias_nstack
Xbias_nstack_0[12] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[12]/vcasc bias_nstack
Xbias_nstack_0[13] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[13]/vcasc bias_nstack
Xbias_nstack_0[14] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[14]/vcasc bias_nstack
Xbias_nstack_0[15] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[15]/vcasc bias_nstack
Xbias_nstack_0[16] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[16]/vcasc bias_nstack
Xbias_nstack_0[17] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[17]/vcasc bias_nstack
Xbias_nstack_0[18] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[18]/vcasc bias_nstack
Xbias_nstack_0[19] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[19]/vcasc bias_nstack
Xbias_nstack_0[20] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[20]/vcasc bias_nstack
Xbias_nstack_0[21] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[21]/vcasc bias_nstack
Xbias_nstack_0[22] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[22]/vcasc bias_nstack
Xbias_nstack_0[23] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[23]/vcasc bias_nstack
Xbias_nstack_0[24] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[24]/vcasc bias_nstack
Xbias_nstack_0[25] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[25]/vcasc bias_nstack
Xbias_nstack_0[26] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[26]/vcasc bias_nstack
Xbias_nstack_0[27] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[27]/vcasc bias_nstack
Xbias_nstack_0[28] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[28]/vcasc bias_nstack
Xbias_nstack_0[29] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[29]/vcasc bias_nstack
Xbias_nstack_0[30] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[30]/vcasc bias_nstack
Xbias_nstack_0[31] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[31]/vcasc bias_nstack
Xbias_nstack_0[32] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[32]/vcasc bias_nstack
Xbias_nstack_0[33] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[33]/vcasc bias_nstack
Xbias_nstack_0[34] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[34]/vcasc bias_nstack
Xbias_nstack_0[35] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[35]/vcasc bias_nstack
Xbias_nstack_0[36] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[36]/vcasc bias_nstack
Xbias_nstack_0[37] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[37]/vcasc bias_nstack
Xbias_nstack_0[38] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[38]/vcasc bias_nstack
Xbias_nstack_0[39] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[39]/vcasc bias_nstack
Xbias_nstack_0[40] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[40]/vcasc bias_nstack
Xbias_nstack_0[41] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[41]/vcasc bias_nstack
Xbias_nstack_0[42] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[42]/vcasc bias_nstack
Xbias_nstack_0[43] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[43]/vcasc bias_nstack
Xbias_nstack_0[44] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[44]/vcasc bias_nstack
Xbias_nstack_0[45] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[45]/vcasc bias_nstack
Xbias_nstack_0[46] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[46]/vcasc bias_nstack
Xbias_nstack_0[47] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[47]/vcasc bias_nstack
Xbias_nstack_0[48] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[48]/vcasc bias_nstack
Xbias_nstack_0[49] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[49]/vcasc bias_nstack
Xbias_nstack_0[50] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[50]/vcasc bias_nstack
Xbias_nstack_0[51] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[51]/vcasc bias_nstack
Xbias_nstack_0[52] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[52]/vcasc bias_nstack
Xbias_nstack_0[53] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[53]/vcasc bias_nstack
Xbias_nstack_0[54] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[54]/vcasc bias_nstack
Xbias_nstack_0[55] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[55]/vcasc bias_nstack
Xbias_nstack_0[56] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[56]/vcasc bias_nstack
Xbias_nstack_0[57] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[57]/vcasc bias_nstack
Xbias_nstack_0[58] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[58]/vcasc bias_nstack
Xbias_nstack_0[59] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[59]/vcasc bias_nstack
Xbias_nstack_0[60] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[60]/vcasc bias_nstack
Xbias_nstack_0[61] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[61]/vcasc bias_nstack
Xbias_nstack_0[62] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[62]/vcasc bias_nstack
Xbias_nstack_0[63] bias_nstack_0[9]/itail ena_bit6 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[63]/vcasc bias_nstack
Xbias_nstack_0[64] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[64]/vcasc bias_nstack
Xbias_nstack_0[65] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[65]/vcasc bias_nstack
Xbias_nstack_0[66] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[66]/vcasc bias_nstack
Xbias_nstack_0[67] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[67]/vcasc bias_nstack
Xbias_nstack_0[68] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[68]/vcasc bias_nstack
Xbias_nstack_0[69] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[69]/vcasc bias_nstack
Xbias_nstack_0[70] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[70]/vcasc bias_nstack
Xbias_nstack_0[71] bias_nstack_0[9]/itail ena_bit3 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[71]/vcasc bias_nstack
Xbias_nstack_0[72] bias_nstack_0[9]/itail ena_bit2 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[72]/vcasc bias_nstack
Xbias_nstack_0[73] bias_nstack_0[9]/itail ena_bit2 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[73]/vcasc bias_nstack
Xbias_nstack_0[74] bias_nstack_0[9]/itail ena_bit2 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[74]/vcasc bias_nstack
Xbias_nstack_0[75] bias_nstack_0[9]/itail ena_bit2 bias_nstack_3[3]/nbias avss_uq2
+ bias_nstack_0[75]/vcasc bias_nstack
Xbias_nstack_1[0] bias_nstack_1[9]/itail avss_uq1 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[0]/vcasc bias_nstack
Xbias_nstack_1[1] bias_nstack_1[9]/itail bias_nstack_1[1]/ena bias_nstack_3[3]/nbias
+ avss_uq1 bias_nstack_1[1]/vcasc bias_nstack
Xbias_nstack_1[2] bias_nstack_1[9]/itail bias_nstack_1[3]/ena bias_nstack_3[3]/nbias
+ avss_uq1 bias_nstack_1[2]/vcasc bias_nstack
Xbias_nstack_1[3] bias_nstack_1[9]/itail bias_nstack_1[3]/ena bias_nstack_3[3]/nbias
+ avss_uq1 bias_nstack_1[3]/vcasc bias_nstack
Xbias_nstack_1[4] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[4]/vcasc bias_nstack
Xbias_nstack_1[5] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[5]/vcasc bias_nstack
Xbias_nstack_1[6] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[6]/vcasc bias_nstack
Xbias_nstack_1[7] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[7]/vcasc bias_nstack
Xbias_nstack_1[8] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[8]/vcasc bias_nstack
Xbias_nstack_1[9] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[9]/vcasc bias_nstack
Xbias_nstack_1[10] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[10]/vcasc bias_nstack
Xbias_nstack_1[11] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[11]/vcasc bias_nstack
Xbias_nstack_1[12] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[12]/vcasc bias_nstack
Xbias_nstack_1[13] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[13]/vcasc bias_nstack
Xbias_nstack_1[14] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[14]/vcasc bias_nstack
Xbias_nstack_1[15] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[15]/vcasc bias_nstack
Xbias_nstack_1[16] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[16]/vcasc bias_nstack
Xbias_nstack_1[17] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[17]/vcasc bias_nstack
Xbias_nstack_1[18] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[18]/vcasc bias_nstack
Xbias_nstack_1[19] bias_nstack_1[9]/itail ena_bit4 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[19]/vcasc bias_nstack
Xbias_nstack_1[20] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[20]/vcasc bias_nstack
Xbias_nstack_1[21] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[21]/vcasc bias_nstack
Xbias_nstack_1[22] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[22]/vcasc bias_nstack
Xbias_nstack_1[23] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[23]/vcasc bias_nstack
Xbias_nstack_1[24] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[24]/vcasc bias_nstack
Xbias_nstack_1[25] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[25]/vcasc bias_nstack
Xbias_nstack_1[26] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[26]/vcasc bias_nstack
Xbias_nstack_1[27] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[27]/vcasc bias_nstack
Xbias_nstack_1[28] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[28]/vcasc bias_nstack
Xbias_nstack_1[29] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[29]/vcasc bias_nstack
Xbias_nstack_1[30] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[30]/vcasc bias_nstack
Xbias_nstack_1[31] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[31]/vcasc bias_nstack
Xbias_nstack_1[32] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[32]/vcasc bias_nstack
Xbias_nstack_1[33] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[33]/vcasc bias_nstack
Xbias_nstack_1[34] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[34]/vcasc bias_nstack
Xbias_nstack_1[35] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[35]/vcasc bias_nstack
Xbias_nstack_1[36] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[36]/vcasc bias_nstack
Xbias_nstack_1[37] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[37]/vcasc bias_nstack
Xbias_nstack_1[38] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[38]/vcasc bias_nstack
Xbias_nstack_1[39] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[39]/vcasc bias_nstack
Xbias_nstack_1[40] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[40]/vcasc bias_nstack
Xbias_nstack_1[41] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[41]/vcasc bias_nstack
Xbias_nstack_1[42] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[42]/vcasc bias_nstack
Xbias_nstack_1[43] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[43]/vcasc bias_nstack
Xbias_nstack_1[44] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[44]/vcasc bias_nstack
Xbias_nstack_1[45] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[45]/vcasc bias_nstack
Xbias_nstack_1[46] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[46]/vcasc bias_nstack
Xbias_nstack_1[47] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[47]/vcasc bias_nstack
Xbias_nstack_1[48] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[48]/vcasc bias_nstack
Xbias_nstack_1[49] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[49]/vcasc bias_nstack
Xbias_nstack_1[50] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[50]/vcasc bias_nstack
Xbias_nstack_1[51] bias_nstack_1[9]/itail ena_bit5 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[51]/vcasc bias_nstack
Xbias_nstack_1[52] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[52]/vcasc bias_nstack
Xbias_nstack_1[53] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[53]/vcasc bias_nstack
Xbias_nstack_1[54] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[54]/vcasc bias_nstack
Xbias_nstack_1[55] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[55]/vcasc bias_nstack
Xbias_nstack_1[56] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[56]/vcasc bias_nstack
Xbias_nstack_1[57] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[57]/vcasc bias_nstack
Xbias_nstack_1[58] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[58]/vcasc bias_nstack
Xbias_nstack_1[59] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[59]/vcasc bias_nstack
Xbias_nstack_1[60] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[60]/vcasc bias_nstack
Xbias_nstack_1[61] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[61]/vcasc bias_nstack
Xbias_nstack_1[62] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[62]/vcasc bias_nstack
Xbias_nstack_1[63] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[63]/vcasc bias_nstack
Xbias_nstack_1[64] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[64]/vcasc bias_nstack
Xbias_nstack_1[65] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[65]/vcasc bias_nstack
Xbias_nstack_1[66] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[66]/vcasc bias_nstack
Xbias_nstack_1[67] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[67]/vcasc bias_nstack
Xbias_nstack_1[68] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[68]/vcasc bias_nstack
Xbias_nstack_1[69] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[69]/vcasc bias_nstack
Xbias_nstack_1[70] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[70]/vcasc bias_nstack
Xbias_nstack_1[71] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[71]/vcasc bias_nstack
Xbias_nstack_1[72] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[72]/vcasc bias_nstack
Xbias_nstack_1[73] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[73]/vcasc bias_nstack
Xbias_nstack_1[74] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[74]/vcasc bias_nstack
Xbias_nstack_1[75] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[75]/vcasc bias_nstack
Xbias_nstack_1[76] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[76]/vcasc bias_nstack
Xbias_nstack_1[77] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[77]/vcasc bias_nstack
Xbias_nstack_1[78] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[78]/vcasc bias_nstack
Xbias_nstack_1[79] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[79]/vcasc bias_nstack
Xbias_nstack_1[80] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[80]/vcasc bias_nstack
Xbias_nstack_1[81] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[81]/vcasc bias_nstack
Xbias_nstack_1[82] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[82]/vcasc bias_nstack
Xbias_nstack_1[83] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[83]/vcasc bias_nstack
Xbias_nstack_1[84] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[84]/vcasc bias_nstack
Xbias_nstack_1[85] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[85]/vcasc bias_nstack
Xbias_nstack_1[86] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[86]/vcasc bias_nstack
Xbias_nstack_1[87] bias_nstack_1[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq1
+ bias_nstack_1[87]/vcasc bias_nstack
Xsky130_fd_sc_hvl__decap_4_8 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xbias_nstack_2[0] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[0]/vcasc
+ bias_nstack
Xbias_nstack_2[1] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[1]/vcasc
+ bias_nstack
Xbias_nstack_2[2] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[2]/vcasc
+ bias_nstack
Xbias_nstack_2[3] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[3]/vcasc
+ bias_nstack
Xbias_nstack_2[4] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[4]/vcasc
+ bias_nstack
Xbias_nstack_2[5] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[5]/vcasc
+ bias_nstack
Xbias_nstack_2[6] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[6]/vcasc
+ bias_nstack
Xbias_nstack_2[7] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[7]/vcasc
+ bias_nstack
Xbias_nstack_2[8] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[8]/vcasc
+ bias_nstack
Xbias_nstack_2[9] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[9]/vcasc
+ bias_nstack
Xbias_nstack_2[10] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[10]/vcasc
+ bias_nstack
Xbias_nstack_2[11] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[11]/vcasc
+ bias_nstack
Xbias_nstack_2[12] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[12]/vcasc
+ bias_nstack
Xbias_nstack_2[13] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[13]/vcasc
+ bias_nstack
Xbias_nstack_2[14] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[14]/vcasc
+ bias_nstack
Xbias_nstack_2[15] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[15]/vcasc
+ bias_nstack
Xbias_nstack_2[16] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[16]/vcasc
+ bias_nstack
Xbias_nstack_2[17] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[17]/vcasc
+ bias_nstack
Xbias_nstack_2[18] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[18]/vcasc
+ bias_nstack
Xbias_nstack_2[19] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[19]/vcasc
+ bias_nstack
Xbias_nstack_2[20] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[20]/vcasc
+ bias_nstack
Xbias_nstack_2[21] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[21]/vcasc
+ bias_nstack
Xbias_nstack_2[22] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[22]/vcasc
+ bias_nstack
Xbias_nstack_2[23] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[23]/vcasc
+ bias_nstack
Xbias_nstack_2[24] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[24]/vcasc
+ bias_nstack
Xbias_nstack_2[25] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[25]/vcasc
+ bias_nstack
Xbias_nstack_2[26] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[26]/vcasc
+ bias_nstack
Xbias_nstack_2[27] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[27]/vcasc
+ bias_nstack
Xbias_nstack_2[28] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[28]/vcasc
+ bias_nstack
Xbias_nstack_2[29] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[29]/vcasc
+ bias_nstack
Xbias_nstack_2[30] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[30]/vcasc
+ bias_nstack
Xbias_nstack_2[31] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[31]/vcasc
+ bias_nstack
Xbias_nstack_2[32] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[32]/vcasc
+ bias_nstack
Xbias_nstack_2[33] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[33]/vcasc
+ bias_nstack
Xbias_nstack_2[34] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[34]/vcasc
+ bias_nstack
Xbias_nstack_2[35] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[35]/vcasc
+ bias_nstack
Xbias_nstack_2[36] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[36]/vcasc
+ bias_nstack
Xbias_nstack_2[37] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[37]/vcasc
+ bias_nstack
Xbias_nstack_2[38] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[38]/vcasc
+ bias_nstack
Xbias_nstack_2[39] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[39]/vcasc
+ bias_nstack
Xbias_nstack_2[40] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[40]/vcasc
+ bias_nstack
Xbias_nstack_2[41] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[41]/vcasc
+ bias_nstack
Xbias_nstack_2[42] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[42]/vcasc
+ bias_nstack
Xbias_nstack_2[43] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[43]/vcasc
+ bias_nstack
Xbias_nstack_2[44] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[44]/vcasc
+ bias_nstack
Xbias_nstack_2[45] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[45]/vcasc
+ bias_nstack
Xbias_nstack_2[46] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[46]/vcasc
+ bias_nstack
Xbias_nstack_2[47] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[47]/vcasc
+ bias_nstack
Xbias_nstack_2[48] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[48]/vcasc
+ bias_nstack
Xbias_nstack_2[49] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[49]/vcasc
+ bias_nstack
Xbias_nstack_2[50] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[50]/vcasc
+ bias_nstack
Xbias_nstack_2[51] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[51]/vcasc
+ bias_nstack
Xbias_nstack_2[52] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[52]/vcasc
+ bias_nstack
Xbias_nstack_2[53] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[53]/vcasc
+ bias_nstack
Xbias_nstack_2[54] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[54]/vcasc
+ bias_nstack
Xbias_nstack_2[55] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[55]/vcasc
+ bias_nstack
Xbias_nstack_2[56] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[56]/vcasc
+ bias_nstack
Xbias_nstack_2[57] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[57]/vcasc
+ bias_nstack
Xbias_nstack_2[58] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[58]/vcasc
+ bias_nstack
Xbias_nstack_2[59] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[59]/vcasc
+ bias_nstack
Xbias_nstack_2[60] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[60]/vcasc
+ bias_nstack
Xbias_nstack_2[61] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[61]/vcasc
+ bias_nstack
Xbias_nstack_2[62] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[62]/vcasc
+ bias_nstack
Xbias_nstack_2[63] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[63]/vcasc
+ bias_nstack
Xbias_nstack_2[64] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[64]/vcasc
+ bias_nstack
Xbias_nstack_2[65] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[65]/vcasc
+ bias_nstack
Xbias_nstack_2[66] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[66]/vcasc
+ bias_nstack
Xbias_nstack_2[67] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[67]/vcasc
+ bias_nstack
Xbias_nstack_2[68] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[68]/vcasc
+ bias_nstack
Xbias_nstack_2[69] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[69]/vcasc
+ bias_nstack
Xbias_nstack_2[70] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[70]/vcasc
+ bias_nstack
Xbias_nstack_2[71] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[71]/vcasc
+ bias_nstack
Xbias_nstack_2[72] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[72]/vcasc
+ bias_nstack
Xbias_nstack_2[73] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[73]/vcasc
+ bias_nstack
Xbias_nstack_2[74] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[74]/vcasc
+ bias_nstack
Xbias_nstack_2[75] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[75]/vcasc
+ bias_nstack
Xbias_nstack_2[76] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[76]/vcasc
+ bias_nstack
Xbias_nstack_2[77] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[77]/vcasc
+ bias_nstack
Xbias_nstack_2[78] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[78]/vcasc
+ bias_nstack
Xbias_nstack_2[79] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[79]/vcasc
+ bias_nstack
Xbias_nstack_2[80] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[80]/vcasc
+ bias_nstack
Xbias_nstack_2[81] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[81]/vcasc
+ bias_nstack
Xbias_nstack_2[82] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[82]/vcasc
+ bias_nstack
Xbias_nstack_2[83] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[83]/vcasc
+ bias_nstack
Xbias_nstack_2[84] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[84]/vcasc
+ bias_nstack
Xbias_nstack_2[85] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[85]/vcasc
+ bias_nstack
Xbias_nstack_2[86] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[86]/vcasc
+ bias_nstack
Xbias_nstack_2[87] bias_nstack_2[9]/itail ena_bit7 bias_nstack_3[3]/nbias avss bias_nstack_2[87]/vcasc
+ bias_nstack
Xsky130_fd_sc_hvl__decap_4_9 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xbias_nstack_3[0] bias_nstack_3[3]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq0
+ bias_nstack_3[0]/vcasc bias_nstack
Xbias_nstack_3[1] bias_nstack_3[3]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq0
+ bias_nstack_3[1]/vcasc bias_nstack
Xbias_nstack_3[2] bias_nstack_3[3]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq0
+ bias_nstack_3[2]/vcasc bias_nstack
Xbias_nstack_3[3] bias_nstack_3[3]/itail ena_bit7 bias_nstack_3[3]/nbias avss_uq0
+ bias_nstack_3[3]/vcasc bias_nstack
Xsky130_fd_sc_hvl__inv_2_0 ena_bit7 dvss dvss avdd_uq2 avdd_uq2 enb_bit7 sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_1 ena_bit3 dvss dvss avdd_uq2 avdd_uq2 enb_bit3 sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|0] ena[7] dvdd dvss avdd_uq2 avdd_uq2 ena_bit7
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|0] ena[6] dvdd dvss avdd_uq2 avdd_uq2 ena_bit6
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[2|0] ena[5] dvdd dvss avdd_uq2 avdd_uq2 ena_bit5
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[3|0] ena[4] dvdd dvss avdd_uq2 avdd_uq2 ena_bit4
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|1] ena[3] dvdd dvss avdd_uq2 avdd_uq2 ena_bit3
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|1] ena[2] dvdd dvss avdd_uq2 avdd_uq2 ena_bit2
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[2|1] ena[1] dvdd dvss avdd_uq2 avdd_uq2 bias_nstack_1[3]/ena
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[3|1] ena[0] dvdd dvss avdd_uq2 avdd_uq2 bias_nstack_1[1]/ena
+ avdd_uq2 dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__inv_2_3 ena_bit5 dvss dvss avdd_uq2 avdd_uq2 enb_bit5 sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_2 ena_bit6 dvss dvss avdd_uq2 avdd_uq2 enb_bit6 sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_4 bias_nstack_1[1]/ena dvss dvss avdd_uq2 avdd_uq2 bias_pstack_1[1]/enb
+ sky130_fd_sc_hvl__inv_2
Xbias_pstack_0[0] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[0]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[1] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[1]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[2] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[2]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[3] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[3]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[4] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[4]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[5] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[5]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[6] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[6]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[7] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[7]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[8] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[8]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[9] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[9]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[10] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[10]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[11] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[11]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[12] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[12]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[13] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[13]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[14] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[14]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[15] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[15]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[16] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[16]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[17] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[17]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[18] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[18]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[19] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[19]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[20] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[20]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[21] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[21]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[22] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[22]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[23] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[23]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[24] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[24]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[25] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[25]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[26] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[26]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[27] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[27]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[28] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[28]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[29] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[29]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[30] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[30]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[31] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[31]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[32] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[32]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[33] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[33]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[34] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[34]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[35] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[35]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[36] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[36]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[37] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[37]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[38] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[38]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[39] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[39]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[40] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[40]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[41] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[41]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[42] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[42]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[43] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[43]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[44] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[44]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[45] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[45]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[46] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[46]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[47] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[47]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[48] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[48]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[49] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[49]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[50] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[50]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[51] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[51]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[52] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[52]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[53] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[53]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[54] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[54]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[55] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[55]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[56] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[56]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[57] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[57]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[58] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[58]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[59] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[59]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[60] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[60]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[61] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[61]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[62] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[62]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[63] bias_pstack_3[3]/pcasc enb_bit6 bias_pstack_0[9]/itail bias_pstack_0[63]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[64] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[64]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[65] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[65]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[66] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[66]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[67] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[67]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[68] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[68]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[69] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[69]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[70] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[70]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[71] bias_pstack_3[3]/pcasc enb_bit3 bias_pstack_0[9]/itail bias_pstack_0[71]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[72] bias_pstack_3[3]/pcasc enb_bit2 bias_pstack_0[9]/itail bias_pstack_0[72]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[73] bias_pstack_3[3]/pcasc enb_bit2 bias_pstack_0[9]/itail bias_pstack_0[73]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[74] bias_pstack_3[3]/pcasc enb_bit2 bias_pstack_0[9]/itail bias_pstack_0[74]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_0[75] bias_pstack_3[3]/pcasc enb_bit2 bias_pstack_0[9]/itail bias_pstack_0[75]/vcasc
+ bias_pstack_3[3]/pbias avss_uq2 avdd_uq2 bias_pstack
Xbias_pstack_1[0] bias_pstack_3[3]/pcasc avdd_uq1 bias_pstack_1[9]/itail bias_pstack_1[0]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[1] bias_pstack_3[3]/pcasc bias_pstack_1[1]/enb bias_pstack_1[9]/itail
+ bias_pstack_1[1]/vcasc bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[2] bias_pstack_3[3]/pcasc bias_pstack_1[3]/enb bias_pstack_1[9]/itail
+ bias_pstack_1[2]/vcasc bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[3] bias_pstack_3[3]/pcasc bias_pstack_1[3]/enb bias_pstack_1[9]/itail
+ bias_pstack_1[3]/vcasc bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[4] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[4]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[5] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[5]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[6] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[6]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[7] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[7]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[8] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[8]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[9] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[9]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[10] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[10]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[11] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[11]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[12] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[12]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[13] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[13]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[14] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[14]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[15] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[15]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[16] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[16]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[17] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[17]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[18] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[18]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[19] bias_pstack_3[3]/pcasc enb_bit4 bias_pstack_1[9]/itail bias_pstack_1[19]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[20] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[20]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[21] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[21]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[22] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[22]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[23] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[23]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[24] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[24]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[25] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[25]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[26] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[26]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[27] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[27]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[28] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[28]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[29] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[29]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[30] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[30]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[31] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[31]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[32] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[32]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[33] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[33]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[34] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[34]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[35] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[35]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[36] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[36]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[37] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[37]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[38] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[38]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[39] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[39]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[40] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[40]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[41] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[41]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[42] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[42]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[43] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[43]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[44] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[44]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[45] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[45]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[46] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[46]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[47] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[47]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[48] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[48]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[49] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[49]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[50] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[50]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[51] bias_pstack_3[3]/pcasc enb_bit5 bias_pstack_1[9]/itail bias_pstack_1[51]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[52] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[52]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[53] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[53]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[54] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[54]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[55] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[55]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[56] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[56]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[57] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[57]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[58] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[58]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[59] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[59]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[60] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[60]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[61] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[61]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[62] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[62]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[63] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[63]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[64] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[64]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[65] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[65]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[66] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[66]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[67] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[67]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[68] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[68]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[69] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[69]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[70] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[70]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[71] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[71]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[72] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[72]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[73] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[73]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[74] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[74]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[75] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[75]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[76] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[76]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[77] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[77]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[78] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[78]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[79] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[79]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[80] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[80]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[81] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[81]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[82] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[82]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[83] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[83]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[84] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[84]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[85] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[85]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[86] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[86]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_1[87] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_1[9]/itail bias_pstack_1[87]/vcasc
+ bias_pstack_3[3]/pbias avss_uq1 avdd_uq1 bias_pstack
Xbias_pstack_2[0] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[0]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[1] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[1]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[2] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[2]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[3] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[3]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[4] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[4]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[5] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[5]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[6] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[6]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[7] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[7]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[8] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[8]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[9] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[9]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[10] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[10]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[11] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[11]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[12] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[12]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[13] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[13]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[14] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[14]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[15] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[15]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[16] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[16]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[17] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[17]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[18] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[18]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[19] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[19]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[20] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[20]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[21] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[21]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[22] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[22]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[23] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[23]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[24] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[24]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[25] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[25]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[26] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[26]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[27] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[27]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[28] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[28]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[29] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[29]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[30] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[30]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[31] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[31]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[32] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[32]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[33] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[33]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[34] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[34]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[35] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[35]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[36] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[36]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[37] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[37]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[38] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[38]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[39] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[39]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[40] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[40]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[41] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[41]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[42] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[42]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[43] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[43]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[44] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[44]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[45] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[45]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[46] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[46]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[47] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[47]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[48] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[48]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[49] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[49]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[50] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[50]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[51] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[51]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[52] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[52]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[53] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[53]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[54] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[54]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[55] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[55]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[56] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[56]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[57] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[57]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[58] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[58]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[59] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[59]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[60] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[60]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[61] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[61]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[62] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[62]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[63] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[63]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[64] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[64]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[65] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[65]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[66] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[66]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[67] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[67]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[68] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[68]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[69] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[69]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[70] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[70]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[71] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[71]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[72] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[72]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[73] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[73]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[74] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[74]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[75] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[75]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[76] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[76]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[77] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[77]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[78] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[78]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[79] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[79]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[80] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[80]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[81] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[81]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[82] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[82]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[83] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[83]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[84] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[84]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[85] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[85]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[86] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[86]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xbias_pstack_2[87] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_2[9]/itail bias_pstack_2[87]/vcasc
+ bias_pstack_3[3]/pbias avss avdd bias_pstack
Xsky130_fd_sc_hvl__inv_2_7 ena_bit2 dvss dvss avdd_uq2 avdd_uq2 enb_bit2 sky130_fd_sc_hvl__inv_2
Xbias_pstack_3[0] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_3[3]/itail bias_pstack_3[0]/vcasc
+ bias_pstack_3[3]/pbias avss_uq0 avdd_uq0 bias_pstack
Xbias_pstack_3[1] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_3[3]/itail bias_pstack_3[1]/vcasc
+ bias_pstack_3[3]/pbias avss_uq0 avdd_uq0 bias_pstack
Xbias_pstack_3[2] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_3[3]/itail bias_pstack_3[2]/vcasc
+ bias_pstack_3[3]/pbias avss_uq0 avdd_uq0 bias_pstack
Xbias_pstack_3[3] bias_pstack_3[3]/pcasc enb_bit7 bias_pstack_3[3]/itail bias_pstack_3[3]/vcasc
+ bias_pstack_3[3]/pbias avss_uq0 avdd_uq0 bias_pstack
Xsky130_fd_sc_hvl__decap_4_10 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_0 ena[3] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_11 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_1 ena[7] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_13 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__decap_4_12 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_2 ena[0] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_3 ena[4] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_4 ena[1] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_16 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_5 ena[5] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_17 dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__inv_2_10 ena_bit4 dvss dvss avdd_uq2 avdd_uq2 enb_bit4 sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_6 ena[2] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_2_11 bias_nstack_1[3]/ena dvss dvss avdd_uq2 avdd_uq2 bias_pstack_1[3]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_7 ena[6] dvss dvss avdd_uq2 avdd_uq2 sky130_fd_sc_hvl__diode_2
.ends

.subckt sky130_ef_ip__idac3v_8bit din[6] din[3] din[2] din[0] din[1] din[5] din[4]
+ din[7] ref_sel_vbg ena vbg src_out ref_in avdd snk_out dvdd dvss avss
Xbias_generator_fe_0 bias_generator_fe_0/snk_test0 bias_generator_fe_0/src_test0 vbg
+ ref_in dvss dvss ref_sel_vbg dvdd dvss bias_generator_fe_0/bias_amp_0/out avdd bias_generator_fe_0/bias_amp_0/nbias
+ ena bias_generator_fe_0/bias_pstack_0[9]/pcasc avss bias_generator_fe
Xbias_generator_idac_be_0 avdd dvdd dvss din[6] din[3] din[2] din[0] din[1] din[5]
+ din[4] din[7] avss avdd avdd avdd dvss dvdd dvss dvdd dvss snk_out bias_generator_fe_0/bias_amp_0/nbias
+ bias_generator_fe_0/bias_pstack_0[9]/pcasc src_out src_out src_out snk_out src_out
+ avss snk_out snk_out avss avss bias_generator_fe_0/bias_amp_0/out bias_generator_idac_be
.ends

.subckt sky130_fd_io__pwrdet_lshv2hv_0_pmos1 a_266_290# a_879_132# a_1191_132# w_0_0#
+ a_266_34# a_1091_34#
X0 a_879_132# a_266_290# w_0_0# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1 a_266_34# a_266_290# w_0_0# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=2.84 as=0.42 ps=2.84 w=0.42 l=1
X2 a_266_290# a_266_34# w_0_0# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=2.84 as=0.42 ps=2.84 w=0.42 l=1
X3 a_1191_132# a_1091_34# w_0_0# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X4 w_0_0# a_266_290# a_879_132# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
.ends

.subckt s8_esd_res250_sub_small a_10_2# a_2142_2#
X0 a_10_2# a_2142_2# sky130_fd_pr__res_generic_po w=2 l=10.07
.ends

.subckt s8_esd_res250only_small rout pad
Xs8_esd_res250_sub_small_0 pad rout s8_esd_res250_sub_small
.ends

.subckt sky130_fd_io__pwrdet_vddd s8_esd_res250only_small_0/rout s8_esd_res250only_small_0/pad
Xs8_esd_res250only_small_0 s8_esd_res250only_small_0/rout s8_esd_res250only_small_0/pad
+ s8_esd_res250only_small
.ends

.subckt sky130_fd_io__pwrdet_vddio s8_esd_res250only_small_0/rout s8_esd_res250only_small_0/pad
Xs8_esd_res250only_small_0 s8_esd_res250only_small_0/rout s8_esd_res250only_small_0/pad
+ s8_esd_res250only_small
.ends

.subckt sky130_fd_io__pwrdet_lshv2hv_0_nmos a_65_173# a_833_141# a_1145_141# a_65_63#
+ a_1245_173# a_365_141# a_2978_173# a_2183_355# a_3086_541#
X0 a_465_173# a_365_141# a_65_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X1 a_1245_173# a_1145_141# a_1089_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X2 a_365_141# a_1145_141# a_65_63# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=1.125 pd=4.5 as=0.105 ps=1.03 w=0.75 l=0.5
X3 a_1089_173# a_833_141# a_65_63# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X4 a_1245_173# a_1145_141# a_1089_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=4.5 pd=9 as=0.42 ps=3.28 w=3 l=0.5
X5 a_65_63# a_65_173# a_2978_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X6 a_65_173# a_365_141# a_465_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X7 a_65_63# a_2183_355# a_1145_141# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=1.125 ps=4.5 w=0.75 l=0.5
X8 a_65_63# a_833_141# a_465_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X9 a_1089_173# a_1145_141# a_1245_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X10 a_65_63# a_3086_541# a_1245_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.8
X11 a_65_63# a_1245_173# a_65_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.63 ps=3.84 w=0.42 l=1
X12 a_465_173# a_365_141# a_65_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=4.5 ps=9 w=3 l=0.5
X13 a_833_141# a_3086_541# a_65_63# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X14 a_1245_173# a_65_173# a_65_63# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.63 pd=3.84 as=0.0588 ps=0.7 w=0.42 l=1
.ends

.subckt sky130_fd_io__pwrdet_lshv2hv_0_pmos2 a_626_66# a_336_n32# w_100_0# a_170_66#
X0 w_100_0# a_336_n32# a_170_66# w_100_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.75 ps=3.5 w=0.75 l=0.5
X1 a_626_66# a_170_66# w_100_0# w_100_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.75 pd=3.5 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt sky130_fd_io__top_pwrdetv2 in1_vddd_hv in2_vddd_hv out3_vddio_hv out1_vddio_hv
+ out2_vddio_hv out2_vddd_hv out1_vddd_hv in1_vddio_hv vddio_present_vddd_hv vddd_present_vddio_hv
+ tie_lo_esd rst_por_hv_n out3_vddd_hv in3_vddio_hv in2_vddio_hv in3_vddd_hv vssio_q
+ vccd vddd1 vssa vddio_q vddd2 vssd
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos1_0 m1_2293_2703# m1_2213_2623# m1_1977_10035#
+ vddio_q a_5004_11122# a_4058_10886# sky130_fd_io__pwrdet_lshv2hv_0_pmos1
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos1_1 m1_771_556# m1_697_476# m1_627_392# vddd1
+ a_6944_17954# a_6025_19417# sky130_fd_io__pwrdet_lshv2hv_0_pmos1
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos1_2 m1_1104_1007# m1_1032_923# m1_957_843# vddd1
+ a_6927_12695# a_6025_19417# sky130_fd_io__pwrdet_lshv2hv_0_pmos1
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos1_3 m1_4935_2408# m1_4577_2542# m1_4264_2542#
+ vddio_q a_6848_10937# a_4058_10886# sky130_fd_io__pwrdet_lshv2hv_0_pmos1
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos1_4 m1_5874_556# m1_5871_11755# m1_6663_392# vddd1
+ a_6397_12079# a_6025_19417# sky130_fd_io__pwrdet_lshv2hv_0_pmos1
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos1_5 m1_5874_2706# m1_6028_8211# m1_6663_2542#
+ vddio_q a_6848_8377# a_4058_10886# sky130_fd_io__pwrdet_lshv2hv_0_pmos1
Xsky130_fd_io__pwrdet_vddd_0 sky130_fd_io__pwrdet_vddd_0/s8_esd_res250only_small_0/rout
+ vddd2 sky130_fd_io__pwrdet_vddd
Xsky130_fd_io__pwrdet_vddio_0 sky130_fd_io__pwrdet_vddio_0/s8_esd_res250only_small_0/rout
+ vddio_q sky130_fd_io__pwrdet_vddio
Xsky130_fd_io__pwrdet_lshv2hv_0_nmos_0 m1_771_556# m1_627_392# m1_1352_1358# vssd
+ a_6944_17954# m1_1408_1468# m1_697_476# in3_vddio_hv a_6025_19417# sky130_fd_io__pwrdet_lshv2hv_0_nmos
Xsky130_fd_io__pwrdet_lshv2hv_0_nmos_1 m1_2293_2703# m1_1977_10035# m2_4976_1949#
+ vssd a_5004_11122# m1_1973_2325# m1_2213_2623# in3_vddd_hv a_4058_10886# sky130_fd_io__pwrdet_lshv2hv_0_nmos
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos2_0 m1_1408_1468# in3_vddio_hv vddio_q m1_1352_1358#
+ sky130_fd_io__pwrdet_lshv2hv_0_pmos2
Xsky130_fd_io__pwrdet_lshv2hv_0_nmos_2 m1_1104_1007# m1_957_843# m1_1520_1880# vssd
+ a_6927_12695# m1_1464_1672# m1_1032_923# in2_vddio_hv a_6025_19417# sky130_fd_io__pwrdet_lshv2hv_0_nmos
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos2_1 m1_1464_1672# in2_vddio_hv vddio_q m1_1520_1880#
+ sky130_fd_io__pwrdet_lshv2hv_0_pmos2
Xsky130_fd_io__pwrdet_lshv2hv_0_nmos_3 m1_4935_2408# m1_4264_2542# m2_5692_1949# vssd
+ a_6848_10937# m1_5621_1800# m1_4577_2542# in2_vddd_hv a_4058_10886# sky130_fd_io__pwrdet_lshv2hv_0_nmos
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos2_2 m1_1973_2325# in3_vddd_hv vddd2 m2_4976_1949#
+ sky130_fd_io__pwrdet_lshv2hv_0_pmos2
Xsky130_fd_io__pwrdet_lshv2hv_0_nmos_4 m1_5874_2706# m1_6663_2542# m2_6408_1949# vssd
+ a_6848_8377# m1_6340_1800# m1_6028_8211# in1_vddd_hv a_4058_10886# sky130_fd_io__pwrdet_lshv2hv_0_nmos
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos2_3 m1_6340_1800# in1_vddd_hv vddd2 m2_6408_1949#
+ sky130_fd_io__pwrdet_lshv2hv_0_pmos2
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos2_4 m1_5621_1800# in2_vddd_hv vddd2 m2_5692_1949#
+ sky130_fd_io__pwrdet_lshv2hv_0_pmos2
Xsky130_fd_io__pwrdet_lshv2hv_0_nmos_5 m1_5874_556# m1_6663_392# m2_3776_1949# vssd
+ a_6397_12079# m1_3708_1800# m1_5871_11755# in1_vddio_hv a_6025_19417# sky130_fd_io__pwrdet_lshv2hv_0_nmos
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos2_5 m1_3708_1800# in1_vddio_hv vddio_q m2_3776_1949#
+ sky130_fd_io__pwrdet_lshv2hv_0_pmos2
X0 vssa a_2722_25404# a_3304_29317# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X1 a_3304_29317# a_2722_25404# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=10.1 ps=14.04 w=5 l=0.5
X2 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=2
X3 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X4 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X5 vddd1 a_5993_18693# vddio_present_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 a_4404_29317# rst_por_hv_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=2.25 ps=6 w=1.5 l=4
X7 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0 ps=0 w=1 l=4
X8 vssa vssa sky130_fd_pr__res_generic_po w=0.33 l=15.635
X9 a_3935_16143# a_2722_25404# vccd vccd sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X10 vccd a_2722_25404# a_3935_16143# vccd sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X11 out3_vddd_hv a_6944_18110# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X12 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0 ps=0 w=3 l=0.5
X13 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X14 a_3935_16143# a_2722_25404# vccd vccd sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=10.5 ps=17 w=7 l=0.5
X15 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X16 vddio_present_vddd_hv a_5993_18693# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X17 out3_vddio_hv a_4985_10940# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X18 vssa a_3164_16015# a_3196_15715# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=1.5 pd=5 as=1.5 ps=5 w=1 l=8
X19 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X20 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0 ps=0 w=3 l=0.5
X21 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X22 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X23 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X24 a_5011_3767# a_4211_3735# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=4
X25 vddd1 a_6944_18110# out3_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X26 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X27 out3_vddd_hv a_6944_18110# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X28 out1_vddd_hv a_6378_12177# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X29 vssd a_6927_12695# a_6817_12995# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X30 vssd a_6848_9735# out2_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X31 vssa a_4211_3735# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X32 vssa a_2722_25404# a_3935_14683# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=4.5 pd=9 as=4.5 ps=9 w=3 l=8
X33 vddd1 a_6378_12177# out1_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X34 a_3304_29317# a_3164_16015# a_4404_29317# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=2.25 pd=6 as=0.21 ps=1.78 w=1.5 l=4
X35 out2_vddd_hv a_6817_12995# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X36 out2_vddd_hv a_6817_12995# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X37 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X38 a_3634_17232# a_3196_15715# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X39 out3_vddd_hv a_6944_18110# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X40 out2_vddio_hv a_6848_9735# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X41 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X42 out1_vddd_hv a_6378_12177# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X43 vddio_q a_3144_11068# a_4058_10886# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.56 as=0.21 ps=1.78 w=1.5 l=0.5
X44 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X45 out1_vddio_hv a_6848_9111# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X46 vssd a_3634_17232# a_6025_19417# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X47 vssd a_6944_17954# a_6944_18110# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X48 vddd_present_vddio_hv a_3122_10886# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X49 a_3144_11068# a_5011_3767# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=2
X50 a_4058_10886# a_3144_11068# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X51 vssd a_6817_12995# out2_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X52 out1_vddio_hv a_6848_9111# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X53 out3_vddio_hv a_4985_10940# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X54 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X55 vddio_q a_3122_10886# vddd_present_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X56 vddd1 a_6927_12695# a_6817_12995# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X57 out2_vddio_hv a_6848_9735# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X58 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0 ps=0 w=1 l=8
X59 a_6025_19417# a_3634_17232# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X60 vddd1 a_6397_12079# a_6378_12177# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X61 a_4404_29317# a_3164_16015# a_3304_29317# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=2.25 ps=6 w=1.5 l=4
X62 vddio_present_vddd_hv a_5993_18693# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X63 vssd a_5993_18693# vddio_present_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X64 vddio_q a_5004_11122# a_4985_10940# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X65 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X66 vddio_q a_3122_10886# vddd_present_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X67 a_3208_7281# a_3039_3259# a_3139_3291# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=4.5 pd=9 as=4.5 ps=9 w=3 l=8
X68 vddd1 a_3634_17232# a_6025_19417# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X69 tie_lo_esd vssd sky130_fd_pr__res_generic_po w=0.5 l=10.2
X70 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.5
X71 vssa a_3935_16143# a_3164_16015# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7.5 pd=13 as=0.7 ps=5.28 w=5 l=0.5
X72 a_2352_39489# a_9590_39549# sky130_fd_pr__res_generic_po w=0.33 l=1.95k
X73 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0 ps=0 w=3 l=0.5
X74 out3_vddd_hv a_6944_18110# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X75 vssd a_4985_10940# out3_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X76 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0 ps=0 w=3 l=0.5
X77 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0 ps=0 w=3 l=0.5
X78 a_5011_3767# a_4211_3735# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=4
X79 vddd1 a_3164_16015# a_3196_15715# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=1.5 pd=5 as=0.14 ps=1.28 w=1 l=8
X80 vddio_present_vddd_hv a_5993_18693# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X81 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0 ps=0 w=3 l=0.5
X82 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0 ps=0 w=3 l=0.5
X83 vddd1 a_6817_12995# out2_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X84 a_3139_3291# a_3039_3259# a_552_39489# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X85 a_6848_9111# a_6848_8377# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X86 out2_vddd_hv a_6817_12995# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X87 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X88 vccd a_2722_25404# a_3935_16143# vccd sky130_fd_pr__pfet_g5v0d10v5 ad=10.5 pd=17 as=0.98 ps=7.28 w=7 l=0.5
X89 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X90 vddd1 a_6944_18110# out3_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X91 vddd1 a_6944_18110# out3_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X92 vssd a_6944_18110# out3_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X93 vddd1 a_6378_12177# out1_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X94 vssd a_6397_12079# a_6378_12177# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X95 vssd a_6848_9111# out1_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X96 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X97 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X98 out3_vddio_hv a_4985_10940# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X99 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X100 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X101 vddio_q a_6848_9111# out1_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X102 vddio_q a_4985_10940# out3_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X103 out2_vddio_hv a_6848_9735# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X104 vddd1 a_6817_12995# out2_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X105 vddd1 a_3196_15715# a_3634_17232# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X106 vssa a_3196_15715# a_3634_17232# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0.105 ps=1.03 w=0.75 l=0.5
X107 vssa a_3039_3259# a_3938_5381# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=4.5 pd=9 as=4.5 ps=9 w=3 l=8
X108 vssd a_6378_12177# out1_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X109 vddd1 a_6944_17954# a_6944_18110# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X110 vddio_q a_6848_9735# out2_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X111 out1_vddd_hv a_6378_12177# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X112 out1_vddd_hv a_6378_12177# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X113 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X114 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X115 vssd a_3144_11068# a_4058_10886# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0.105 ps=1.03 w=0.75 l=0.5
X116 a_6025_19417# a_3634_17232# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X117 out2_vddd_hv a_6817_12995# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X118 a_4058_10886# a_3144_11068# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X119 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X120 vssa a_4211_3735# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X121 a_3634_17232# a_3196_15715# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X122 vddio_q a_6848_9111# out1_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X123 vddio_q a_4211_3735# a_5011_3767# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=4
X124 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X125 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X126 vssa a_4211_3735# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X127 vddd2 vddd2 vssd sky130_fd_pr__res_generic_nd__hv w=0.3 l=68.84
X128 vssa a_4211_3735# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X129 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0 ps=0 w=0.75 l=0.5
X130 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0 ps=0 w=1.5 l=0.5
X131 vddio_q a_5011_3767# a_3144_11068# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=2
X132 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0 ps=0 w=0.75 l=0.5
X133 vssd a_6378_12177# out1_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X134 vssa a_4211_3735# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X135 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0 ps=0 w=0.75 l=0.5
X136 a_3304_29317# rst_por_hv_n vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=1.5 pd=5 as=1.5 ps=5 w=1 l=1
X137 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X138 out1_vddd_hv a_6378_12177# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X139 vssd a_3144_11068# a_4058_10886# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X140 a_3164_16015# a_3935_16143# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X141 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0 ps=0 w=1.5 l=0.5
X142 vssd a_3122_10886# vddd_present_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X143 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0 ps=0 w=3 l=0.5
X144 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0 ps=0 w=3 l=0.5
X145 vddd1 a_3634_17232# a_5993_18693# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.42 ps=3.56 w=1.5 l=0.5
X146 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0 ps=0 w=1.5 l=0.5
X147 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X148 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0 ps=0 w=3 l=0.5
X149 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0 ps=0 w=0.75 l=0.5
X150 a_552_39489# a_3039_3259# a_3139_3291# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X151 out3_vddd_hv a_6944_18110# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X152 a_3139_3291# a_3039_3259# a_552_39489# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=10.395 ps=16.97 w=7 l=0.5
X153 out2_vddio_hv a_6848_9735# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X154 vddd1 a_6378_12177# out1_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X155 out2_vddio_hv a_6848_9735# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X156 vssd a_3634_17232# a_6025_19417# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0.105 ps=1.03 w=0.75 l=0.5
X157 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X158 out3_vddio_hv a_4985_10940# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X159 vssd a_6848_9735# out2_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X160 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X161 out1_vddio_hv a_6848_9111# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X162 out1_vddio_hv a_6848_9111# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X163 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.5
X164 a_3164_16015# a_3935_16143# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X165 a_9590_39549# vddio_q vssd sky130_fd_pr__res_generic_nd__hv w=0.3 l=1.33932k
X166 a_3304_29317# a_2722_25404# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X167 vddio_q a_6848_9735# out2_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X168 a_3208_7281# a_3039_3259# a_3938_5381# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=4.5 pd=9 as=4.5 ps=9 w=3 l=8
X169 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=2
X170 vssa a_3935_16143# a_3164_16015# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X171 out1_vddd_hv a_6378_12177# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X172 out2_vddio_hv a_6848_9735# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X173 a_4058_10886# a_3144_11068# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X174 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0 ps=0 w=1 l=4
X175 vddd1 a_6378_12177# out1_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X176 vddio_q a_4985_10940# out3_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X177 out2_vddd_hv a_6817_12995# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X178 out2_vddd_hv a_6817_12995# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X179 vddio_q a_6848_8377# a_6848_9111# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X180 vssa a_3304_29317# a_3164_16015# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=2.25 pd=6 as=0.21 ps=1.78 w=1.5 l=4
X181 a_3935_16143# a_2722_25404# vccd vccd sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X182 a_3634_17232# a_3196_15715# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21 ps=2.06 w=0.75 l=0.5
X183 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X184 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X185 vccd a_2722_25404# a_3935_16143# vccd sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X186 vddd1 a_3634_17232# a_6025_19417# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.56 as=0.21 ps=1.78 w=1.5 l=0.5
X187 out3_vddd_hv a_6944_18110# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X188 vddio_q a_3144_11068# a_4058_10886# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X189 vddd_present_vddio_hv a_3122_10886# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X190 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X191 vssd a_5993_18693# vddio_present_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X192 out1_vddio_hv a_6848_9111# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X193 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X194 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X195 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X196 vssd a_6817_12995# out2_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X197 vddio_present_vddd_hv a_5993_18693# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X198 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X199 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X200 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.56 as=0 ps=0 w=1.5 l=0.5
X201 vssd a_3122_10886# vddd_present_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X202 a_6025_19417# a_3634_17232# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X203 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0 ps=0 w=1.5 l=0.5
X204 vddd_present_vddio_hv a_3122_10886# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X205 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0 ps=0 w=3 l=0.5
X206 vddd1 a_3164_16015# a_3304_29317# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.63 pd=3.84 as=0.63 ps=3.84 w=0.42 l=20
X207 vssd a_3634_17232# a_5993_18693# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21 ps=2.06 w=0.75 l=0.5
X208 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X209 a_3164_16015# a_3304_29317# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=2.25 ps=6 w=1.5 l=4
X210 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0 ps=0 w=3 l=0.5
X211 vssd a_6944_18110# out3_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X212 a_552_39489# a_3039_3259# a_3139_3291# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=10.5 pd=17 as=0.98 ps=7.28 w=7 l=0.5
X213 vssd a_5004_11122# a_4985_10940# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X214 a_5835_15413# a_2722_25404# a_3935_16143# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=4.5 pd=9 as=4.5 ps=9 w=3 l=8
X215 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0 ps=0 w=3 l=0.5
X216 a_3935_16143# a_2722_25404# vccd vccd sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X217 vddd1 a_5993_18693# vddio_present_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X218 vddio_q a_4985_10940# out3_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X219 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X220 vssd a_4985_10940# out3_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X221 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X222 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.56 as=0 ps=0 w=1.5 l=0.5
X223 vddio_q a_6848_9111# out1_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X224 a_5835_15413# a_2722_25404# a_3935_14683# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=4.5 pd=9 as=4.5 ps=9 w=3 l=8
X225 a_4211_3735# a_3139_3291# a_3967_4161# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=1.5 pd=5 as=1.5 ps=5 w=1 l=8
X226 out3_vddio_hv a_4985_10940# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X227 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X228 a_3039_3259# sky130_fd_io__pwrdet_vddd_0/s8_esd_res250only_small_0/rout vssd sky130_fd_pr__res_generic_nd__hv w=0.3 l=68.84
X229 vddio_q a_6848_9735# out2_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X230 vddio_q a_6848_9735# out2_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X231 out3_vddio_hv a_4985_10940# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X232 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X233 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0 ps=0 w=1.5 l=0.5
X234 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X235 vddio_q a_4985_10940# out3_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X236 vssa a_5011_3767# a_3144_11068# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=2
X237 vddd1 a_3304_29317# a_3164_16015# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.63 pd=3.84 as=0.63 ps=3.84 w=0.42 l=20
X238 vssa a_2722_25404# a_3304_29317# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X239 vddd1 a_6817_12995# out2_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X240 out1_vddio_hv a_6848_9111# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X241 vddd_present_vddio_hv a_3122_10886# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X242 vssa a_3196_15715# a_3634_17232# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X243 vssd a_3144_11068# a_3122_10886# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21 ps=2.06 w=0.75 l=0.5
X244 a_3196_15715# a_3164_16015# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=1.5 ps=5 w=1 l=8
X245 vddd1 a_6944_18110# out3_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X246 a_6848_9735# a_6848_10937# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X247 vssd a_6848_9111# out1_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X248 a_4211_3735# a_3139_3291# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7.7 pd=16.2 as=7.7 ps=16.2 w=7 l=0.5
X249 vssa rst_por_hv_n a_4404_29317# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=2.25 pd=6 as=0.21 ps=1.78 w=1.5 l=4
X250 vddio_q a_6848_9111# out1_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X251 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X252 vccd a_2722_25404# a_3935_16143# vccd sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X253 vddd1 a_6817_12995# out2_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X254 a_552_39489# a_2352_39489# vssd sky130_fd_pr__res_generic_nd__hv w=0.3 l=3.14938k
X255 vddd1 a_3196_15715# a_3634_17232# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X256 vddio_q a_6848_10937# a_6848_9735# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X257 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X258 a_6025_19417# a_3634_17232# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X259 a_4058_10886# a_3144_11068# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X260 vddio_q a_3144_11068# a_3122_10886# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.42 ps=3.56 w=1.5 l=0.5
X261 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X262 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X263 a_2722_25404# sky130_fd_io__pwrdet_vddio_0/s8_esd_res250only_small_0/rout vssd sky130_fd_pr__res_generic_nd__hv w=0.3 l=277.39001
X264 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X265 a_3634_17232# a_3196_15715# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X266 vddio_q a_3139_3291# a_3967_4161# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=1.5 pd=5 as=1.5 ps=5 w=1 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PXF6AN a_1235_n100# a_n287_n188# a_761_n100#
+ a_819_n188# a_n1077_n188# a_n29_n100# a_345_n188# a_n919_n188# a_977_n188# a_n445_n188#
+ a_n187_n100# a_n1235_n188# a_503_n188# a_n819_n100# a_n603_n188# a_n345_n100# a_1135_n188#
+ a_661_n188# a_n977_n100# a_n1135_n100# a_n761_n188# a_129_n100# a_n503_n100# a_n1293_n100#
+ a_n661_n100# a_287_n100# a_919_n100# a_445_n100# a_1077_n100# a_29_n188# a_n1427_n322#
+ a_n129_n188# a_603_n100# a_187_n188#
X0 a_445_n100# a_345_n188# a_287_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_603_n100# a_503_n188# a_445_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n977_n100# a_n1077_n188# a_n1135_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_n1135_n100# a_n1235_n188# a_n1293_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X4 a_n661_n100# a_n761_n188# a_n819_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_129_n100# a_29_n188# a_n29_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_n187_n100# a_n287_n188# a_n345_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 a_n819_n100# a_n919_n188# a_n977_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 a_n345_n100# a_n445_n188# a_n503_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X9 a_n503_n100# a_n603_n188# a_n661_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X10 a_n29_n100# a_n129_n188# a_n187_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 a_1077_n100# a_977_n188# a_919_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X12 a_761_n100# a_661_n188# a_603_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X13 a_287_n100# a_187_n188# a_129_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X14 a_1235_n100# a_1135_n188# a_1077_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X15 a_919_n100# a_819_n188# a_761_n100# a_n1427_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X5 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12495 pd=1.175 as=0.2184 ps=2.2 w=0.84 l=0.15
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.12495 ps=1.175 w=0.42 l=0.15
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12285 ps=1.17 w=0.84 l=0.15
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1404 pd=1.6 as=0.1137 ps=1.01 w=0.54 l=0.15
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1137 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.10783 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.07438 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12228 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07438 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.12228 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08937 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08937 ps=0.925 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
X0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.09588 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.09588 ps=0.945 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.11213 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.11213 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.27995 ps=1.615 w=1 l=0.15
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.17515 ps=1.265 w=0.65 l=0.15
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.07455 ps=0.775 w=0.42 l=0.15
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X12 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X13 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19627 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.19627 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.10187 ps=0.99 w=0.65 l=0.15
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.1113 ps=1.37 w=0.42 l=0.15
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt brownout_dig VPWR brout_filt dcomp ena force_dis_rc_osc force_ena_rc_osc force_short_oneshot
+ osc_ck otrip[0] otrip[1] otrip[2] vtrip[0] vtrip[1] vtrip[2] osc_ena otrip_decoded[0]
+ otrip_decoded[1] otrip_decoded[3] otrip_decoded[4] otrip_decoded[5] otrip_decoded[6]
+ otrip_decoded[7] outb_unbuf timed_out vtrip_decoded[0] vtrip_decoded[1] vtrip_decoded[2]
+ vtrip_decoded[3] vtrip_decoded[4] vtrip_decoded[5] vtrip_decoded[6] vtrip_decoded[7]
+ otrip_decoded[2] VGND
XFILLER_0_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_062_ net9 net7 net8 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__and3_1
X_045_ net1 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
X_114_ clknet_1_1__leaf_osc_ck _010_ net3 VGND VGND VPWR VPWR cnt\[8\] sky130_fd_sc_hd__dfstp_1
Xoutput31 net31 VGND VGND VPWR VPWR vtrip_decoded[7] sky130_fd_sc_hd__clkbuf_4
Xoutput20 net20 VGND VGND VPWR VPWR otrip_decoded[6] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_044_ net4 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__inv_2
X_061_ net7 net8 net9 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__and3b_1
X_113_ clknet_1_1__leaf_osc_ck _009_ net33 VGND VGND VPWR VPWR cnt\[7\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput21 net21 VGND VGND VPWR VPWR otrip_decoded[7] sky130_fd_sc_hd__buf_2
XFILLER_0_13_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_060_ net8 net7 net9 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__and3b_1
X_043_ net32 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__inv_2
X_112_ clknet_1_0__leaf_osc_ck _008_ net33 VGND VGND VPWR VPWR cnt\[6\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput22 net22 VGND VGND VPWR VPWR outb_unbuf sky130_fd_sc_hd__buf_2
XFILLER_0_13_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_111_ clknet_1_0__leaf_osc_ck _007_ net33 VGND VGND VPWR VPWR cnt\[5\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_12_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput23 net23 VGND VGND VPWR VPWR timed_out sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_15_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_110_ clknet_1_0__leaf_osc_ck _006_ net33 VGND VGND VPWR VPWR cnt\[4\] sky130_fd_sc_hd__dfstp_1
Xoutput24 net24 VGND VGND VPWR VPWR vtrip_decoded[0] sky130_fd_sc_hd__clkbuf_4
Xoutput13 net13 VGND VGND VPWR VPWR osc_ena sky130_fd_sc_hd__buf_2
XFILLER_0_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput25 net25 VGND VGND VPWR VPWR vtrip_decoded[1] sky130_fd_sc_hd__clkbuf_4
Xoutput14 net14 VGND VGND VPWR VPWR otrip_decoded[0] sky130_fd_sc_hd__buf_2
X_099_ cnt\[9\] _022_ cnt\[10\] VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput26 net26 VGND VGND VPWR VPWR vtrip_decoded[2] sky130_fd_sc_hd__clkbuf_4
Xoutput15 net15 VGND VGND VPWR VPWR otrip_decoded[1] sky130_fd_sc_hd__buf_2
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_119__35 VGND VGND VPWR VPWR net35 _119__35/LO sky130_fd_sc_hd__conb_1
X_098_ net23 _023_ _028_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_7_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput27 net27 VGND VGND VPWR VPWR vtrip_decoded[3] sky130_fd_sc_hd__clkbuf_4
Xoutput16 net16 VGND VGND VPWR VPWR otrip_decoded[2] sky130_fd_sc_hd__buf_2
X_097_ cnt\[9\] _022_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__xor2_1
Xoutput28 net28 VGND VGND VPWR VPWR vtrip_decoded[4] sky130_fd_sc_hd__clkbuf_4
Xoutput17 net17 VGND VGND VPWR VPWR otrip_decoded[3] sky130_fd_sc_hd__buf_2
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_096_ cnt\[8\] _035_ net6 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_079_ cnt\[2\] _030_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput29 net29 VGND VGND VPWR VPWR vtrip_decoded[5] sky130_fd_sc_hd__clkbuf_4
Xoutput18 net18 VGND VGND VPWR VPWR otrip_decoded[4] sky130_fd_sc_hd__buf_2
X_095_ _038_ _021_ net38 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_078_ _038_ _040_ net32 VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__a21oi_1
Xoutput19 net19 VGND VGND VPWR VPWR otrip_decoded[5] sky130_fd_sc_hd__buf_2
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout32 clr_cnt VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
X_094_ cnt\[8\] _035_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__xnor2_1
X_077_ _030_ _039_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_11_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_093_ _038_ _020_ net32 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__a21oi_1
Xfanout33 net3 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_4
Xinput1 brout_filt VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_076_ cnt\[1\] cnt\[0\] VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_50 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_059_ net7 net8 net9 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__nor3b_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_092_ cnt\[7\] _034_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__xor2_1
Xinput2 dcomp VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_075_ net39 _038_ net32 VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__a21oi_1
X_058_ net9 net7 net8 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__and3b_1
XFILLER_0_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_074_ net6 net23 VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__nor2_2
X_091_ _038_ _019_ net32 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__a21oi_1
Xinput3 ena VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
X_057_ net9 net7 net8 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__nor3b_1
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_109_ clknet_1_0__leaf_osc_ck _005_ net33 VGND VGND VPWR VPWR cnt\[3\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_090_ _034_ _018_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 force_dis_rc_osc VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_056_ net9 net8 net7 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__nor3b_1
X_073_ net2 net33 VGND VGND VPWR VPWR dcomp_ena_rsb sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_6_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_108_ clknet_1_1__leaf_osc_ck _004_ net33 VGND VGND VPWR VPWR cnt\[2\] sky130_fd_sc_hd__dfstp_1
X_072_ net33 _029_ _037_ net5 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__a31o_1
Xinput5 force_ena_rc_osc VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_055_ net9 net7 net8 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__nor3_1
X_107_ clknet_1_0__leaf_osc_ck _003_ net33 VGND VGND VPWR VPWR cnt\[1\] sky130_fd_sc_hd__dfstp_1
X_118__34 VGND VGND VPWR VPWR _118__34/HI net34 sky130_fd_sc_hd__conb_1
Xinput6 force_short_oneshot VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
X_071_ dcomp_retimed net2 net23 VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_054_ dcomp_retimed net23 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__and2b_1
X_106_ clknet_1_0__leaf_osc_ck _002_ net33 VGND VGND VPWR VPWR cnt\[0\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_070_ net12 net11 net10 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__and3_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 otrip[0] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
X_053_ cnt\[8\] cnt\[11\] _035_ _036_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__and4_2
XFILLER_0_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput10 vtrip[0] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dlymetal6s2s_1
X_105_ net1 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_1_1__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
Xinput8 otrip[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
X_052_ cnt\[9\] cnt\[10\] VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__and2_1
X_104_ net23 _026_ _027_ _028_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__o31a_1
X_121_ clknet_1_1__leaf_osc_ck net2 dcomp_ena_rsb VGND VGND VPWR VPWR dcomp_retimed
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput11 vtrip[1] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput9 otrip[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
X_051_ cnt\[4\] cnt\[7\] _031_ _033_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__and4_1
X_120_ clknet_1_0__leaf_osc_ck net37 _001_ VGND VGND VPWR VPWR clr_cnt_sb sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 vtrip[2] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlymetal6s2s_1
X_103_ _036_ _022_ cnt\[11\] VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 clr_cnt_sb VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
X_050_ _032_ _033_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__nand2_1
X_102_ cnt\[11\] _036_ _022_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__and3b_1
Xclkbuf_0_osc_ck osc_ck VGND VGND VPWR VPWR clknet_0_osc_ck sky130_fd_sc_hd__clkbuf_16
Xhold2 clr_cnt_sb_stg1 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_101_ _028_ net23 _024_ _025_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3 clr_cnt VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_2_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_100_ _036_ _022_ net32 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_5_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold4 cnt\[0\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_089_ cnt\[5\] cnt\[4\] _031_ cnt\[6\] VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_088_ _038_ _017_ net32 VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_9_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_087_ cnt\[5\] _032_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_0__f_osc_ck clknet_0_osc_ck VGND VGND VPWR VPWR clknet_1_0__leaf_osc_ck
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_086_ _038_ _016_ net32 VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__a21oi_1
X_069_ net10 net11 net12 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_085_ _032_ _015_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__or2_1
X_068_ net11 net10 net12 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__and3b_1
X_067_ net11 net10 net12 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__nor3b_1
X_084_ cnt\[4\] _031_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_13_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_119_ clknet_1_0__leaf_osc_ck net35 _000_ VGND VGND VPWR VPWR clr_cnt_sb_stg1 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_083_ _038_ _014_ net32 VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_049_ cnt\[5\] cnt\[6\] VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__and2_1
X_066_ net12 net11 net10 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__and3b_1
X_118_ clknet_1_0__leaf_osc_ck net34 net36 VGND VGND VPWR VPWR clr_cnt sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_4_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_065_ net12 net10 net11 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__nor3b_1
X_082_ _031_ _042_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_048_ cnt\[4\] _031_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__and2_1
X_117_ clknet_1_1__leaf_osc_ck _013_ net3 VGND VGND VPWR VPWR cnt\[11\] sky130_fd_sc_hd__dfstp_1
X_081_ cnt\[1\] cnt\[0\] cnt\[2\] cnt\[3\] VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_064_ net12 net11 net10 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__nor3b_1
X_047_ cnt\[1\] cnt\[0\] cnt\[3\] cnt\[2\] VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__and4_1
X_116_ clknet_1_1__leaf_osc_ck _012_ net3 VGND VGND VPWR VPWR cnt\[10\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_063_ net12 net11 net10 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__nor3_1
X_080_ _038_ _041_ net32 VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_046_ cnt\[1\] cnt\[0\] VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__nand2_1
X_115_ clknet_1_1__leaf_osc_ck _011_ net3 VGND VGND VPWR VPWR cnt\[9\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput30 net30 VGND VGND VPWR VPWR vtrip_decoded[6] sky130_fd_sc_hd__clkbuf_4
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_V6EN4F a_n321_n322# a_n29_n100# a_n187_n100#
+ a_129_n100# a_29_n188# a_n129_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n188# a_n187_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_XTZQRT a_n287_n188# a_761_n100# a_n29_n100# a_345_n188#
+ a_n953_n322# a_n445_n188# a_n187_n100# a_503_n188# a_n819_n100# a_n603_n188# a_n345_n100#
+ a_661_n188# a_n761_n188# a_129_n100# a_n503_n100# a_n661_n100# a_287_n100# a_445_n100#
+ a_29_n188# a_n129_n188# a_603_n100# a_187_n188#
X0 a_445_n100# a_345_n188# a_287_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_603_n100# a_503_n188# a_445_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n661_n100# a_n761_n188# a_n819_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_129_n100# a_29_n188# a_n29_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_n187_n100# a_n287_n188# a_n345_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_n345_n100# a_n445_n188# a_n503_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_n503_n100# a_n603_n188# a_n661_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 a_n29_n100# a_n129_n188# a_n187_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 a_761_n100# a_661_n188# a_603_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X9 a_287_n100# a_187_n188# a_129_n100# a_n953_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A LVPWR VGND VPB VPWR X VPWR_uq0 VGND_uq0 VNB
X0 a_30_1337# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X1 VGND_uq0 a_30_1337# a_30_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.17887 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X2 VGND_uq0 a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X3 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X4 VGND_uq0 a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X5 VGND_uq0 a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X6 VGND A a_30_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.17887 pd=1.26 as=0.1197 ps=1.41 w=0.42 l=0.5
X7 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X8 a_389_141# a_30_207# VGND_uq0 VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.17887 ps=1.26 w=0.75 l=0.5
X9 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X10 LVPWR a_389_141# X LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1568 pd=1.4 as=0.2968 ps=2.77 w=1.12 l=0.15
X11 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.17887 ps=1.26 w=0.75 l=0.5
X12 VGND_uq0 a_389_141# X VNB sky130_fd_pr__nfet_01v8 ad=0.1961 pd=2.01 as=0.1961 ps=2.01 w=0.74 l=0.15
X13 LVPWR a_389_1337# a_389_141# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.2968 ps=2.77 w=1.12 l=0.15
X14 a_30_207# a_30_1337# VPWR_uq0 VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1197 ps=1.41 w=0.42 l=0.5
X15 a_389_1337# a_389_141# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2968 pd=2.77 as=0.1568 ps=1.4 w=1.12 l=0.15
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_K8JYEQ a_n3678_n531# a_296_n557# a_950_n531#
+ a_n2374_n557# a_3976_n531# a_2908_n531# a_n1306_n557# a_n3442_n557# a_n2076_n531#
+ a_n3144_n531# a_2610_n557# a_1542_n557# a_n950_n557# a_n1008_n531# a_n4212_n531#
+ a_3442_n531# a_2374_n531# a_1306_n531# a_n652_n531# a_1898_n557# a_n3798_n557# a_2966_n557#
+ a_772_n531# a_118_n557# a_3798_n531# a_n1720_n531# a_n1128_n557# a_n2196_n557# a_n3264_n557#
+ a_1364_n557# a_3500_n557# a_2432_n557# a_n772_n557# a_2196_n531# a_n474_n531# a_n4034_n531#
+ a_3264_n531# a_1128_n531# a_830_n557# a_3856_n557# a_2788_n557# a_n1840_n557# a_594_n531#
+ a_n1542_n531# a_n2610_n531# a_n3086_n557# a_2254_n557# a_1186_n557# a_n594_n557#
+ a_n2018_n557# a_n4154_n557# a_1840_n531# a_3322_n557# a_3086_n531# a_n296_n531#
+ a_n1898_n531# a_n2966_n531# a_4154_n531# a_2018_n531# a_60_n531# a_652_n557# a_3678_n557#
+ a_n1662_n557# a_n2730_n557# a_n1364_n531# a_n60_n557# a_416_n531# a_n2432_n531#
+ a_1662_n531# a_n3500_n531# a_3144_n557# a_2076_n557# a_1008_n557# a_2730_n531# a_n416_n557#
+ a_n2788_n531# a_n3856_n531# a_474_n557# a_n118_n531# a_n1484_n557# a_n2552_n557#
+ a_n3620_n557# a_238_n531# a_n1186_n531# a_n2254_n531# a_1720_n557# a_n3322_n531#
+ a_n4346_n691# a_2552_n531# a_1484_n531# a_n830_n531# a_4034_n557# a_n3976_n557#
+ a_3620_n531# a_n238_n557# a_n2908_n557#
X0 a_n3856_n531# a_n3976_n557# a_n4034_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 a_n2610_n531# a_n2730_n557# a_n2788_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_n2254_n531# a_n2374_n557# a_n2432_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X3 a_2196_n531# a_2076_n557# a_2018_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X4 a_n652_n531# a_n772_n557# a_n830_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X5 a_2018_n531# a_1898_n557# a_1840_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 a_n1008_n531# a_n1128_n557# a_n1186_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X7 a_594_n531# a_474_n557# a_416_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_3264_n531# a_3144_n557# a_3086_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X9 a_n3322_n531# a_n3442_n557# a_n3500_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X10 a_60_n531# a_n60_n557# a_n118_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X11 a_3086_n531# a_2966_n557# a_2908_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X12 a_1484_n531# a_1364_n557# a_1306_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X13 a_n1542_n531# a_n1662_n557# a_n1720_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X14 a_2552_n531# a_2432_n557# a_2374_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X15 a_950_n531# a_830_n557# a_772_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X16 a_3620_n531# a_3500_n557# a_3442_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X17 a_n3678_n531# a_n3798_n557# a_n3856_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X18 a_n830_n531# a_n950_n557# a_n1008_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X19 a_n2076_n531# a_n2196_n557# a_n2254_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X20 a_n474_n531# a_n594_n557# a_n652_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X21 a_1840_n531# a_1720_n557# a_1662_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X22 a_416_n531# a_296_n557# a_238_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X23 a_n3500_n531# a_n3620_n557# a_n3678_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X24 a_n3144_n531# a_n3264_n557# a_n3322_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X25 a_2908_n531# a_2788_n557# a_2730_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X26 a_4154_n531# a_4034_n557# a_3976_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X27 a_n1898_n531# a_n2018_n557# a_n2076_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X28 a_n296_n531# a_n416_n557# a_n474_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X29 a_1306_n531# a_1186_n557# a_1128_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X30 a_n1720_n531# a_n1840_n557# a_n1898_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X31 a_n1364_n531# a_n1484_n557# a_n1542_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X32 a_238_n531# a_118_n557# a_60_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X33 a_3976_n531# a_3856_n557# a_3798_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X34 a_n2788_n531# a_n2908_n557# a_n2966_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X35 a_n2432_n531# a_n2552_n557# a_n2610_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X36 a_2374_n531# a_2254_n557# a_2196_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X37 a_1128_n531# a_1008_n557# a_950_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X38 a_n1186_n531# a_n1306_n557# a_n1364_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X39 a_772_n531# a_652_n557# a_594_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X40 a_3442_n531# a_3322_n557# a_3264_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X41 a_1662_n531# a_1542_n557# a_1484_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X42 a_n2966_n531# a_n3086_n557# a_n3144_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X43 a_2730_n531# a_2610_n557# a_2552_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X44 a_n4034_n531# a_n4154_n557# a_n4212_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X45 a_n118_n531# a_n238_n557# a_n296_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X46 a_3798_n531# a_3678_n557# a_3620_n531# a_n4346_n691# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_4Z8MHY a_652_n562# a_n1186_n536# a_238_n536#
+ a_n1662_n562# a_3678_n562# a_n2254_n536# a_n2730_n562# a_n3322_n536# a_n60_n562#
+ a_1484_n536# a_2552_n536# a_n830_n536# a_3620_n536# w_n4412_n762# a_2076_n562# a_3144_n562#
+ a_1008_n562# a_n3678_n536# a_n416_n562# a_950_n536# a_474_n562# a_3976_n536# a_2908_n536#
+ a_n1484_n562# a_n2076_n536# a_n2552_n562# a_n3144_n536# a_n1008_n536# a_n3620_n562#
+ a_n4212_n536# a_1720_n562# a_2374_n536# a_n652_n536# a_1306_n536# a_3442_n536# a_n3976_n562#
+ a_4034_n562# a_n238_n562# a_772_n536# a_n2908_n562# a_296_n562# a_3798_n536# a_n1720_n536#
+ a_n2374_n562# a_n3442_n562# a_n1306_n562# a_n4034_n536# a_1542_n562# a_2196_n536#
+ a_n474_n536# a_2610_n562# a_n950_n562# a_1128_n536# a_3264_n536# a_n3798_n562# a_594_n536#
+ a_1898_n562# a_2966_n562# a_n1542_n536# a_n2610_n536# a_118_n562# a_n2196_n562#
+ a_1840_n536# a_n3264_n562# a_n1128_n562# a_1364_n562# a_n1898_n536# a_n296_n536#
+ a_2432_n562# a_n2966_n536# a_n772_n562# a_3086_n536# a_3500_n562# a_2018_n536# a_4154_n536#
+ a_60_n536# a_830_n562# a_2788_n562# a_n1364_n536# a_416_n536# a_n1840_n562# a_3856_n562#
+ a_n2432_n536# a_n3500_n536# a_1662_n536# a_n3086_n562# a_2730_n536# a_n4154_n562#
+ a_n2018_n562# a_1186_n562# a_2254_n562# a_n2788_n536# a_n594_n562# a_3322_n562#
+ a_n3856_n536# a_n118_n536#
X0 a_2552_n536# a_2432_n562# a_2374_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 a_3620_n536# a_3500_n562# a_3442_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_n3678_n536# a_n3798_n562# a_n3856_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X3 a_950_n536# a_830_n562# a_772_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X4 a_n830_n536# a_n950_n562# a_n1008_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X5 a_n2076_n536# a_n2196_n562# a_n2254_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 a_n474_n536# a_n594_n562# a_n652_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X7 a_1840_n536# a_1720_n562# a_1662_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_n3500_n536# a_n3620_n562# a_n3678_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X9 a_n3144_n536# a_n3264_n562# a_n3322_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X10 a_416_n536# a_296_n562# a_238_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X11 a_2908_n536# a_2788_n562# a_2730_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X12 a_n1898_n536# a_n2018_n562# a_n2076_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X13 a_n296_n536# a_n416_n562# a_n474_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X14 a_1306_n536# a_1186_n562# a_1128_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X15 a_4154_n536# a_4034_n562# a_3976_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X16 a_n1720_n536# a_n1840_n562# a_n1898_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X17 a_n1364_n536# a_n1484_n562# a_n1542_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X18 a_3976_n536# a_3856_n562# a_3798_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X19 a_238_n536# a_118_n562# a_60_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X20 a_n2788_n536# a_n2908_n562# a_n2966_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X21 a_2374_n536# a_2254_n562# a_2196_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X22 a_n2432_n536# a_n2552_n562# a_n2610_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X23 a_1128_n536# a_1008_n562# a_950_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X24 a_n1186_n536# a_n1306_n562# a_n1364_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X25 a_3442_n536# a_3322_n562# a_3264_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X26 a_772_n536# a_652_n562# a_594_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X27 a_1662_n536# a_1542_n562# a_1484_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X28 a_n2966_n536# a_n3086_n562# a_n3144_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X29 a_2730_n536# a_2610_n562# a_2552_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X30 a_n118_n536# a_n238_n562# a_n296_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X31 a_n4034_n536# a_n4154_n562# a_n4212_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X32 a_3798_n536# a_3678_n562# a_3620_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X33 a_n3856_n536# a_n3976_n562# a_n4034_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X34 a_n2610_n536# a_n2730_n562# a_n2788_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X35 a_2196_n536# a_2076_n562# a_2018_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X36 a_n2254_n536# a_n2374_n562# a_n2432_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X37 a_n652_n536# a_n772_n562# a_n830_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X38 a_2018_n536# a_1898_n562# a_1840_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X39 a_n1008_n536# a_n1128_n562# a_n1186_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X40 a_3264_n536# a_3144_n562# a_3086_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X41 a_n3322_n536# a_n3442_n562# a_n3500_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X42 a_60_n536# a_n60_n562# a_n118_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X43 a_594_n536# a_474_n562# a_416_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X44 a_3086_n536# a_2966_n562# a_2908_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X45 a_1484_n536# a_1364_n562# a_1306_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X46 a_n1542_n536# a_n1662_n562# a_n1720_n536# w_n4412_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_WY4TLZ a_n919_n536# a_207_n562# a_n1217_n562#
+ w_n1653_n762# a_n385_n536# a_1039_n536# a_n861_n562# a_n1453_n536# a_505_n536# a_1275_n562#
+ a_29_n562# a_n1039_n562# a_n683_n562# a_n207_n536# a_741_n562# a_327_n536# a_n1275_n536#
+ a_1097_n562# a_n505_n562# a_n29_n536# a_n1097_n536# a_563_n562# a_149_n536# a_1395_n536#
+ a_n741_n536# a_919_n562# a_861_n536# a_n327_n562# a_385_n562# a_n1395_n562# a_1217_n536#
+ a_n563_n536# a_683_n536# a_n149_n562#
X0 a_n1275_n536# a_n1395_n562# a_n1453_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X1 a_n741_n536# a_n861_n562# a_n919_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_n1097_n536# a_n1217_n562# a_n1275_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X3 a_1039_n536# a_919_n562# a_861_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X4 a_683_n536# a_563_n562# a_505_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X5 a_n29_n536# a_n149_n562# a_n207_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 a_n563_n536# a_n683_n562# a_n741_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X7 a_n919_n536# a_n1039_n562# a_n1097_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_505_n536# a_385_n562# a_327_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X9 a_n385_n536# a_n505_n562# a_n563_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X10 a_1395_n536# a_1275_n562# a_1217_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X11 a_327_n536# a_207_n562# a_149_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X12 a_149_n536# a_29_n562# a_n29_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X13 a_861_n536# a_741_n562# a_683_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X14 a_n207_n536# a_n327_n562# a_n385_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X15 a_1217_n536# a_1097_n562# a_1039_n536# w_n1653_n762# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_9VZRJ2 a_n7134_n3916# a_n8646_3484# a_7230_3484#
+ a_n5244_3484# a_8364_n3916# a_12144_3484# a_n7512_n3916# a_6096_n3916# a_n9024_3484#
+ a_n5244_n3916# a_n12048_n3916# a_8742_n3916# a_6474_n3916# a_n330_n3916# a_n708_n3916#
+ a_n12426_n3916# a_48_n3916# a_n5622_n3916# a_n7890_3484# a_7986_3484# a_n12804_3484#
+ a_4584_3484# a_n2598_3484# a_n3354_n3916# a_n10158_n3916# a_n13182_3484# a_1182_3484#
+ a_6852_n3916# a_n12804_n3916# a_11388_n3916# a_4584_n3916# a_n1086_n3916# a_8364_3484#
+ a_n10536_n3916# a_n3732_n3916# a_n6378_3484# a_11766_n3916# a_4962_n3916# a_n1464_n3916#
+ a_n10914_n3916# a_2694_n3916# a_n1842_n3916# a_n9780_n3916# a_n1842_3484# a_1938_3484#
+ a_48_3484# a_n10536_3484# a_n5622_3484# a_5718_3484# a_9498_3484# a_n2220_3484#
+ a_n7890_n3916# a_2316_3484# a_6096_3484# a_12522_3484# a_9120_n3916# a_n9402_3484#
+ a_n6000_3484# a_n6000_n3916# a_7230_n3916# a_7608_n3916# a_426_n3916# a_4962_3484#
+ a_1560_3484# a_n2976_3484# a_804_n3916# a_n4110_n3916# a_8742_3484# a_n6756_3484#
+ a_5340_3484# a_12144_n3916# a_n3354_3484# a_5340_n3916# a_5718_n3916# a_n13312_n4046#
+ a_n12048_3484# a_10254_3484# a_3072_n3916# a_9120_3484# a_12522_n3916# a_n2220_n3916#
+ a_n7134_3484# a_426_3484# a_10254_n3916# a_3450_n3916# a_3828_n3916# a_12900_n3916#
+ a_n708_3484# a_1182_n3916# a_n8268_n3916# a_10632_n3916# a_n10914_3484# a_2694_3484#
+ a_n11292_3484# a_9498_n3916# a_n8646_n3916# a_n9780_3484# a_1560_n3916# a_1938_n3916#
+ a_9876_3484# a_6474_3484# a_12900_3484# a_n4488_3484# a_3072_3484# a_9876_n3916#
+ a_n1086_3484# a_n6378_n3916# a_11388_3484# a_n8268_3484# a_n13182_n3916# a_n6756_n3916#
+ a_n330_3484# a_7986_n3916# a_n4488_n3916# a_n11292_n3916# a_n4866_n3916# a_n2598_n3916#
+ a_n3732_3484# a_3828_3484# a_n11670_n3916# a_n12426_3484# a_10632_3484# a_n2976_n3916#
+ a_n7512_3484# a_7608_3484# a_804_3484# a_n4110_3484# a_4206_3484# a_4206_n3916#
+ a_11010_3484# a_11010_n3916# a_n11670_3484# a_2316_n3916# a_n9024_n3916# a_6852_3484#
+ a_3450_3484# a_n4866_3484# a_n9402_n3916# a_n1464_3484# a_n10158_3484# a_11766_3484#
X0 a_n9024_3484# a_n9024_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X1 a_9876_3484# a_9876_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X2 a_6474_3484# a_6474_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X3 a_n11670_3484# a_n11670_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X4 a_n7890_3484# a_n7890_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X5 a_n330_3484# a_n330_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X6 a_3072_3484# a_3072_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X7 a_5718_3484# a_5718_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X8 a_8742_3484# a_8742_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X9 a_n11292_3484# a_n11292_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X10 a_n10536_3484# a_n10536_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X11 a_n4488_3484# a_n4488_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X12 a_2316_3484# a_2316_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X13 a_5340_3484# a_5340_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X14 a_12144_3484# a_12144_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X15 a_n12804_3484# a_n12804_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X16 a_n6756_3484# a_n6756_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X17 a_n1086_3484# a_n1086_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X18 a_n5622_3484# a_n5622_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X19 a_n3354_3484# a_n3354_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X20 a_11010_3484# a_11010_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X21 a_9498_3484# a_9498_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X22 a_6096_3484# a_6096_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X23 a_7608_3484# a_7608_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X24 a_8364_3484# a_8364_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X25 a_n13182_3484# a_n13182_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X26 a_n10158_3484# a_n10158_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X27 a_n9780_3484# a_n9780_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X28 a_4206_3484# a_4206_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X29 a_7230_3484# a_7230_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X30 a_n12426_3484# a_n12426_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X31 a_n8646_3484# a_n8646_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X32 a_n6378_3484# a_n6378_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X33 a_n7512_3484# a_n7512_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X34 a_n5244_3484# a_n5244_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X35 a_n2220_3484# a_n2220_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X36 a_1938_3484# a_1938_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X37 a_2694_3484# a_2694_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X38 a_4962_3484# a_4962_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X39 a_1560_3484# a_1560_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X40 a_11766_3484# a_11766_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X41 a_n2976_3484# a_n2976_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X42 a_48_3484# a_48_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X43 a_10632_3484# a_10632_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X44 a_n1842_3484# a_n1842_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X45 a_12900_3484# a_12900_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X46 a_804_3484# a_804_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X47 a_9120_3484# a_9120_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X48 a_n12048_3484# a_n12048_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X49 a_n8268_3484# a_n8268_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X50 a_n9402_3484# a_n9402_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X51 a_n7134_3484# a_n7134_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X52 a_n4110_3484# a_n4110_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X53 a_7986_3484# a_7986_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X54 a_4584_3484# a_4584_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X55 a_6852_3484# a_6852_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X56 a_n6000_3484# a_n6000_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X57 a_n708_3484# a_n708_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X58 a_1182_3484# a_1182_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X59 a_3450_3484# a_3450_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X60 a_3828_3484# a_3828_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X61 a_11388_3484# a_11388_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X62 a_n10914_3484# a_n10914_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X63 a_n4866_3484# a_n4866_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X64 a_n2598_3484# a_n2598_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X65 a_10254_3484# a_10254_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X66 a_n1464_3484# a_n1464_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X67 a_12522_3484# a_12522_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X68 a_n3732_3484# a_n3732_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X69 a_426_3484# a_426_n3916# a_n13312_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z__0 a_100_n100# a_n292_n322# a_n158_n100#
+ a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n292_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt rstring_mux vout_brout ena otrip_decoded_avdd[7] otrip_decoded_avdd[6] otrip_decoded_avdd[5]
+ otrip_decoded_avdd[4] otrip_decoded_avdd[3] otrip_decoded_avdd[2] otrip_decoded_avdd[1]
+ vtrip_decoded_avdd[7] vtrip_decoded_avdd[6] vtrip_decoded_avdd[5] vtrip_decoded_avdd[4]
+ vtrip_decoded_avdd[3] vtrip_decoded_avdd[2] vtrip_decoded_avdd[1] vtrip_decoded_avdd[0]
+ vout_vunder vtop otrip_decoded_avdd[0] avdd avss
Xsky130_fd_pr__nfet_g5v0d10v5_K8JYEQ_0 vout_brout vtrip_decoded_avdd[0] vout_vunder
+ otrip_decoded_avdd[3] vtrip7 vtrip5 otrip_decoded_avdd[5] otrip_decoded_avdd[1]
+ vout_brout vout_brout avss avss otrip_decoded_avdd[6] vout_brout vout_brout vtrip6
+ vtrip4 vtrip2 vout_brout vtrip_decoded_avdd[3] avss vtrip_decoded_avdd[5] vtrip1
+ vtrip_decoded_avdd[0] vout_vunder vout_brout avss avss avss vtrip_decoded_avdd[2]
+ vtrip_decoded_avdd[6] vtrip_decoded_avdd[4] otrip_decoded_avdd[6] vout_vunder vout_brout
+ vtrip0 vout_vunder vout_vunder vtrip_decoded_avdd[1] vtrip_decoded_avdd[7] vtrip_decoded_avdd[5]
+ otrip_decoded_avdd[4] vout_vunder vout_brout vout_brout otrip_decoded_avdd[2] vtrip_decoded_avdd[4]
+ vtrip_decoded_avdd[2] avss otrip_decoded_avdd[4] otrip_decoded_avdd[0] vtrip3 vtrip_decoded_avdd[6]
+ vout_vunder vtrip7 vtrip4 vtrip2 vout_vunder vout_vunder vout_vunder vtrip_decoded_avdd[1]
+ avss avss avss vtrip5 avss vout_vunder vtrip3 vout_vunder vtrip1 avss avss avss
+ vout_vunder otrip_decoded_avdd[7] vout_brout vout_brout avss vout_brout otrip_decoded_avdd[5]
+ otrip_decoded_avdd[3] otrip_decoded_avdd[1] vtrip0 vout_brout vout_brout vtrip_decoded_avdd[3]
+ vout_brout avss vout_vunder vout_vunder vtrip6 vtrip_decoded_avdd[7] otrip_decoded_avdd[0]
+ vout_vunder otrip_decoded_avdd[7] otrip_decoded_avdd[2] sky130_fd_pr__nfet_g5v0d10v5_K8JYEQ
Xsky130_fd_pr__pfet_g5v0d10v5_4Z8MHY_0 vtrip_decoded_b_avdd[1] vout_brout vtrip0 avdd
+ avdd vout_brout avdd vout_brout avdd vout_vunder vout_vunder vtrip6 vout_vunder
+ avdd avdd avdd avdd vout_brout otrip_decoded_b_avdd[7] vout_vunder avdd vtrip7 vtrip5
+ otrip_decoded_b_avdd[5] vout_brout otrip_decoded_b_avdd[3] vout_brout vout_brout
+ otrip_decoded_b_avdd[1] vout_brout vtrip_decoded_b_avdd[3] vtrip4 vout_brout vtrip2
+ vtrip6 otrip_decoded_b_avdd[0] vtrip_decoded_b_avdd[7] otrip_decoded_b_avdd[7] vtrip1
+ otrip_decoded_b_avdd[2] vtrip_decoded_b_avdd[0] vout_vunder vout_brout otrip_decoded_b_avdd[3]
+ otrip_decoded_b_avdd[1] otrip_decoded_b_avdd[5] vtrip0 avdd vout_vunder vout_brout
+ avdd otrip_decoded_b_avdd[6] vout_vunder vout_vunder avdd vout_vunder vtrip_decoded_b_avdd[3]
+ vtrip_decoded_b_avdd[5] vout_brout vout_brout vtrip_decoded_b_avdd[0] avdd vtrip3
+ avdd avdd vtrip_decoded_b_avdd[2] vtrip4 vtrip7 vtrip_decoded_b_avdd[4] vtrip2 otrip_decoded_b_avdd[6]
+ vout_vunder vtrip_decoded_b_avdd[6] vout_vunder vout_vunder vout_vunder vtrip_decoded_b_avdd[1]
+ vtrip_decoded_b_avdd[5] vtrip5 vout_vunder otrip_decoded_b_avdd[4] vtrip_decoded_b_avdd[7]
+ vtrip3 vtrip1 vout_vunder otrip_decoded_b_avdd[2] vout_vunder otrip_decoded_b_avdd[0]
+ otrip_decoded_b_avdd[4] vtrip_decoded_b_avdd[2] vtrip_decoded_b_avdd[4] vout_brout
+ avdd vtrip_decoded_b_avdd[6] vout_brout vout_brout sky130_fd_pr__pfet_g5v0d10v5_4Z8MHY
Xsky130_fd_pr__pfet_g5v0d10v5_WY4TLZ_0 vtop ena_b ena_b avdd avdd avdd ena_b avdd
+ vtop ena_b ena_b ena_b ena_b vtop ena_b avdd vtop ena_b ena_b avdd avdd ena_b vtop
+ avdd avdd ena_b vtop ena_b ena_b ena_b vtop vtop avdd ena_b sky130_fd_pr__pfet_g5v0d10v5_WY4TLZ
Xsky130_fd_sc_hvl__inv_1_0[0] otrip_decoded_avdd[0] avss avss avdd avdd otrip_decoded_b_avdd[0]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[1] otrip_decoded_avdd[1] avss avss avdd avdd otrip_decoded_b_avdd[1]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[2] otrip_decoded_avdd[2] avss avss avdd avdd otrip_decoded_b_avdd[2]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[3] otrip_decoded_avdd[3] avss avss avdd avdd otrip_decoded_b_avdd[3]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[4] otrip_decoded_avdd[4] avss avss avdd avdd otrip_decoded_b_avdd[4]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[5] otrip_decoded_avdd[5] avss avss avdd avdd otrip_decoded_b_avdd[5]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[6] otrip_decoded_avdd[6] avss avss avdd avdd otrip_decoded_b_avdd[6]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[7] otrip_decoded_avdd[7] avss avss avdd avdd otrip_decoded_b_avdd[7]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[8] vtrip_decoded_avdd[0] avss avss avdd avdd vtrip_decoded_b_avdd[0]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[9] vtrip_decoded_avdd[1] avss avss avdd avdd vtrip_decoded_b_avdd[1]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[10] vtrip_decoded_avdd[2] avss avss avdd avdd vtrip_decoded_b_avdd[2]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[11] vtrip_decoded_avdd[3] avss avss avdd avdd vtrip_decoded_b_avdd[3]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[12] vtrip_decoded_avdd[4] avss avss avdd avdd vtrip_decoded_b_avdd[4]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[13] vtrip_decoded_avdd[5] avss avss avdd avdd vtrip_decoded_b_avdd[5]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[14] vtrip_decoded_avdd[6] avss avss avdd avdd vtrip_decoded_b_avdd[6]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_0[15] vtrip_decoded_avdd[7] avss avss avdd avdd vtrip_decoded_b_avdd[7]
+ sky130_fd_sc_hvl__inv_1
Xsky130_fd_sc_hvl__inv_1_1 ena avss avss avdd avdd ena_b sky130_fd_sc_hvl__inv_1
Xsky130_fd_pr__res_xhigh_po_1p41_9VZRJ2_0 m1_6950_n3340# m1_5060_4059# m1_20936_4059#
+ m1_8840_4059# m1_22070_n3340# m1_26228_4059# m1_6194_n3340# m1_19802_n3340# m1_5060_4059#
+ m1_8462_n3340# m1_1658_n3340# m1_22826_n3340# m1_20558_n3340# vtrip0 m1_12998_n3340#
+ m1_1658_n3340# vtrip0 m1_8462_n3340# m1_5816_4059# m1_21692_4059# m1_1280_4059#
+ m1_18668_4059# m1_11108_4059# m1_10730_n3340# m1_3926_n3340# vtop vtrip3 m1_20558_n3340#
+ m1_902_n3340# m1_25094_n3340# m1_18290_n3340# m1_12998_n3340# m1_22448_4059# m1_3170_n3340#
+ m1_9974_n3340# m1_7328_4059# m1_25850_n3340# m1_19046_n3340# m1_12242_n3340# m1_3170_n3340#
+ m1_16778_n3340# m1_12242_n3340# m1_3926_n3340# m1_11864_4059# vtrip5 vtrip1 m1_3548_4059#
+ m1_8084_4059# m1_19424_4059# m1_23204_4059# m1_11864_4059# m1_6194_n3340# vtrip7
+ m1_20180_4059# m1_26228_4059# m1_22826_n3340# m1_4304_4059# m1_8084_4059# m1_7706_n3340#
+ m1_21314_n3340# m1_21314_n3340# vtrip2 m1_18668_4059# vtrip5 m1_11108_4059# vtrip2
+ m1_9974_n3340# m1_22448_4059# m1_7328_4059# m1_19424_4059# m1_25850_n3340# m1_10352_4059#
+ m1_19046_n3340# m1_19802_n3340# avss m1_2036_4059# m1_23960_4059# m1_16778_n3340#
+ m1_23204_4059# m1_26606_n3340# m1_11486_n3340# m1_6572_4059# vtrip1 m1_24338_n3340#
+ m1_17534_n3340# m1_17534_n3340# m1_26606_n3340# m1_13376_4059# vtrip4 m1_5438_n3340#
+ m1_24338_n3340# m1_2792_4059# vtrip7 m1_2792_4059# m1_23582_n3340# m1_5438_n3340#
+ m1_4304_4059# vtrip4 vtrip6 m1_23960_4059# m1_20180_4059# avss m1_9596_4059# m1_17156_4059#
+ m1_23582_n3340# m1_12620_4059# m1_7706_n3340# m1_25472_4059# m1_5816_4059# m1_902_n3340#
+ m1_6950_n3340# m1_13376_4059# m1_22070_n3340# m1_9218_n3340# m1_2414_n3340# m1_9218_n3340#
+ m1_11486_n3340# m1_10352_4059# m1_17912_4059# m1_2414_n3340# m1_1280_4059# m1_24716_4059#
+ m1_10730_n3340# m1_6572_4059# m1_21692_4059# vtrip3 m1_9596_4059# m1_17912_4059#
+ m1_18290_n3340# m1_24716_4059# m1_25094_n3340# m1_2036_4059# vtrip6 m1_4682_n3340#
+ m1_20936_4059# m1_17156_4059# m1_8840_4059# m1_4682_n3340# m1_12620_4059# m1_3548_4059#
+ m1_25472_4059# sky130_fd_pr__res_xhigh_po_1p41_9VZRJ2
Xsky130_fd_pr__nfet_g5v0d10v5_CD9S2Z_0 avss avss vtop ena_b sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z__0
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_SCV3UK a_50_n131# a_n50_n157# a_n526_n243# a_n108_n131#
+ a_n266_n131# a_n424_n131# a_208_n131# a_108_n157# a_n208_n157# a_366_n131# a_266_n157#
+ a_n366_n157#
X0 a_n108_n131# a_n208_n157# a_n266_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_208_n131# a_108_n157# a_50_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n266_n131# a_n366_n157# a_n424_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_366_n131# a_266_n157# a_208_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X4 a_50_n131# a_n50_n157# a_n108_n131# a_n526_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_BZXTE7 a_208_n64# a_n108_n64# a_998_n64# a_n898_n64#
+ a_108_n161# a_50_n64# a_n208_n161# a_266_n161# a_n424_n64# a_524_n64# a_898_n161#
+ a_n366_n161# a_424_n161# a_n998_n161# a_n266_n64# a_366_n64# a_n524_n161# a_582_n161#
+ a_n50_n161# a_840_n64# a_n740_n64# a_n682_n161# a_740_n161# a_682_n64# a_n582_n64#
+ a_n840_n161# w_n1194_n284# a_n1056_n64#
X0 a_n898_n64# a_n998_n161# a_n1056_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X1 a_n582_n64# a_n682_n161# a_n740_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_50_n64# a_n50_n161# a_n108_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_n740_n64# a_n840_n161# a_n898_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_n266_n64# a_n366_n161# a_n424_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_n424_n64# a_n524_n161# a_n582_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_n108_n64# a_n208_n161# a_n266_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 a_998_n64# a_898_n161# a_840_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X8 a_682_n64# a_582_n161# a_524_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X9 a_840_n64# a_740_n161# a_682_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X10 a_366_n64# a_266_n161# a_208_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 a_524_n64# a_424_n161# a_366_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X12 a_208_n64# a_108_n161# a_50_n64# w_n1194_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt schmitt_trigger in out dvdd dvss
Xsky130_fd_pr__nfet_01v8_SCV3UK_1 m out dvss dvss m dvss dvss dvss in out m in sky130_fd_pr__nfet_01v8_SCV3UK
Xsky130_fd_pr__pfet_01v8_BZXTE7_0 dvdd dvdd out m out m in out dvdd dvdd m in dvdd
+ in m m in m out dvdd dvdd in m out m in dvdd dvdd sky130_fd_pr__pfet_01v8_BZXTE7
.ends

.subckt sky130_fd_pr__pfet_01v8_MA8JJJ a_18_n136# a_n33_95# w_n112_n198# a_n76_n136#
X0 a_18_n136# a_n33_95# a_n76_n136# w_n112_n198# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.18
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_V6VPPZ a_n1842_n10916# a_n708_n10916# a_426_10484#
+ a_804_10484# a_n1464_n10916# a_n1972_n11046# a_1182_10484# a_n1086_n10916# a_1560_10484#
+ a_48_n10916# a_804_n10916# a_n330_10484# a_n708_10484# a_1560_n10916# a_48_10484#
+ a_426_n10916# a_n1086_10484# a_n1464_10484# a_1182_n10916# a_n1842_10484# a_n330_n10916#
X0 a_426_10484# a_426_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X1 a_n708_10484# a_n708_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X2 a_1560_10484# a_1560_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X3 a_n1086_10484# a_n1086_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X4 a_n1842_10484# a_n1842_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X5 a_n330_10484# a_n330_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X6 a_1182_10484# a_1182_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X7 a_48_10484# a_48_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X8 a_804_10484# a_804_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
X9 a_n1464_10484# a_n1464_n10916# a_n1972_n11046# sky130_fd_pr__res_xhigh_po_1p41 l=105
.ends

.subckt sky130_fd_pr__pfet_01v8_LAUYMQ w_n161_n200# a_n125_n100# a_66_n100# a_15_131#
+ a_n30_n100# a_n81_n197#
X0 a_n30_n100# a_n81_n197# a_n125_n100# w_n161_n200# sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.295 ps=2.59 w=1 l=0.18
X1 a_66_n100# a_15_131# a_n30_n100# w_n161_n200# sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.15 ps=1.3 w=1 l=0.18
.ends

.subckt sky130_fd_pr__pfet_01v8_C64SS5 a_287_n64# a_n187_n64# a_129_n64# w_n539_n164#
+ a_29_n161# a_n129_n161# a_187_n161# a_n29_n64# a_n287_n161# a_n503_n64# a_345_n161#
+ a_n345_n64# a_445_n64# a_n445_n161#
X0 a_129_n64# a_29_n161# a_n29_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n187_n64# a_n287_n161# a_n345_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n345_n64# a_n445_n161# a_n503_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_n29_n64# a_n129_n161# a_n187_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_287_n64# a_187_n161# a_129_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_445_n64# a_345_n161# a_287_n64# w_n539_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_LUWKLG c2_n3269_n19000# m4_n3349_n19080#
X0 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X1 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X2 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X3 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X4 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
X5 c2_n3269_n19000# m4_n3349_n19080# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
.ends

.subckt sky130_fd_pr__pfet_01v8_2XUZHN a_n73_n100# w_n109_n162# a_15_n100# a_n15_n126#
X0 a_15_n100# a_n15_n126# a_n73_n100# w_n109_n162# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_C68ZY6 a_208_n64# a_n108_n64# a_108_n161# w_n618_n164#
+ a_50_n64# a_n208_n161# a_266_n161# a_n424_n64# a_524_n64# a_n366_n161# a_424_n161#
+ a_n266_n64# a_366_n64# a_n524_n161# a_n50_n161# a_n582_n64#
X0 a_50_n64# a_n50_n161# a_n108_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n266_n64# a_n366_n161# a_n424_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n424_n64# a_n524_n161# a_n582_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_n108_n64# a_n208_n161# a_n266_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_366_n64# a_266_n161# a_208_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_524_n64# a_424_n161# a_366_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X6 a_208_n64# a_108_n161# a_50_n64# w_n618_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_C6GQGA w_n154_n164# a_n118_n64# a_60_n64# a_n60_n161#
X0 a_60_n64# a_n60_n161# a_n118_n64# w_n154_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.6
.ends

.subckt sky130_fd_pr__pfet_01v8_9QCJ55 a_358_n64# a_n158_n64# a_158_n161# a_n358_n161#
+ a_n100_n161# w_n452_n164# a_100_n64# a_n416_n64#
X0 a_100_n64# a_n100_n161# a_n158_n64# w_n452_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X1 a_358_n64# a_158_n161# a_100_n64# w_n452_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X2 a_n158_n64# a_n358_n161# a_n416_n64# w_n452_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_MLERZ7 a_50_n136# a_n108_n136# a_n50_n162# w_n144_n198#
X0 a_50_n136# a_n50_n162# a_n108_n136# w_n144_n198# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt rc_osc dvdd out ena dvss
Xsky130_fd_pr__pfet_01v8_MA8JJJ_0 dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_MA8JJJ
Xsky130_fd_pr__res_xhigh_po_1p41_V6VPPZ_0 vr m1_2270_n4# m1_23669_n1138# m1_23669_n1138#
+ m1_2270_752# dvss m1_23669_n1894# m1_2270_752# m1_23669_n1894# m1_2270_n760# m1_2270_n1516#
+ m1_23669_n382# m1_23669_374# in m1_23669_n382# m1_2270_n760# m1_23669_374# m1_23669_1130#
+ m1_2270_n1516# m1_23669_1130# m1_2270_n4# sky130_fd_pr__res_xhigh_po_1p41_V6VPPZ
Xsky130_fd_pr__pfet_01v8_LAUYMQ_0 dvdd dvdd vr ena_b out dvdd sky130_fd_pr__pfet_01v8_LAUYMQ
Xsky130_fd_pr__pfet_01v8_C64SS5_0 m dvdd dvdd dvdd in in in m in dvdd in m dvdd in
+ sky130_fd_pr__pfet_01v8_C64SS5
Xsky130_fd_pr__cap_mim_m3_2_LUWKLG_0 in dvss sky130_fd_pr__cap_mim_m3_2_LUWKLG
Xsky130_fd_pr__pfet_01v8_2XUZHN_0 in dvdd dvdd ena sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_C68ZY6_0 out n n dvdd dvdd m n n out m n dvdd dvdd dvdd m
+ m sky130_fd_pr__pfet_01v8_C68ZY6
Xsky130_fd_pr__pfet_01v8_C6GQGA_0 dvdd dvdd ena_b ena sky130_fd_pr__pfet_01v8_C6GQGA
Xsky130_fd_pr__pfet_01v8_9QCJ55_0 m m n n n dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_9QCJ55
Xsky130_fd_pr__pfet_01v8_MLERZ7_0 vr ena_b dvdd dvdd sky130_fd_pr__pfet_01v8_MLERZ7
X0 dvss dvss m dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 m n dvss dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X2 dvss ena ena_b dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X3 out ena vr dvss sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.1475 ps=1.295 w=1 l=0.18
X4 dvss dvss n dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 dvss in m dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 n m dvss dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 dvss dvss out dvss sky130_fd_pr__nfet_01v8 ad=0.1475 pd=1.295 as=0.15 ps=1.3 w=1 l=0.18
X8 m in dvss dvss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.1475 ps=1.295 w=1 l=0.5
X9 vr dvss dvss dvss sky130_fd_pr__nfet_01v8 ad=0.1475 pd=1.295 as=0.145 ps=1.29 w=1 l=0.6
X10 out n dvss dvss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_DVQADA a_48_n3916# a_n330_n3916# a_n708_n3916#
+ a_1182_3484# a_n2598_3484# a_n3354_n3916# a_n1086_n3916# a_n3732_n3916# a_n1464_n3916#
+ a_2694_n3916# a_n1842_n3916# a_n3862_n4046# a_1938_3484# a_48_3484# a_n1842_3484#
+ a_n2220_3484# a_2316_3484# a_426_n3916# a_1560_3484# a_n2976_3484# a_804_n3916#
+ a_n3354_3484# a_3072_n3916# a_426_3484# a_n2220_n3916# a_3450_n3916# a_n708_3484#
+ a_2694_3484# a_1182_n3916# a_1938_n3916# a_1560_n3916# a_3072_3484# a_n1086_3484#
+ a_n330_3484# a_n2598_n3916# a_n3732_3484# a_804_3484# a_n2976_n3916# a_2316_n3916#
+ a_3450_3484# a_n1464_3484#
X0 a_n330_3484# a_n330_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X1 a_3072_3484# a_3072_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X2 a_2316_3484# a_2316_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X3 a_n1086_3484# a_n1086_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X4 a_n3354_3484# a_n3354_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X5 a_n2220_3484# a_n2220_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X6 a_1938_3484# a_1938_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X7 a_2694_3484# a_2694_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X8 a_1560_3484# a_1560_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X9 a_n2976_3484# a_n2976_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X10 a_48_3484# a_48_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X11 a_n1842_3484# a_n1842_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X12 a_804_3484# a_804_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X13 a_n708_3484# a_n708_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X14 a_1182_3484# a_1182_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X15 a_3450_3484# a_3450_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X16 a_n2598_3484# a_n2598_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X17 a_n1464_3484# a_n1464_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X18 a_n3732_3484# a_n3732_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
X19 a_426_3484# a_426_n3916# a_n3862_n4046# sky130_fd_pr__res_xhigh_po_1p41 l=35
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_XZ4X25 a_n887_n588# a_n429_n588# a_487_n588#
+ a_n945_n500# a_29_n588# a_n487_n500# a_n1079_n722# a_n29_n500# a_887_n500# a_429_n500#
X0 a_n29_n500# a_n429_n588# a_n487_n500# a_n1079_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X1 a_429_n500# a_29_n588# a_n29_n500# a_n1079_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X2 a_887_n500# a_487_n588# a_429_n500# a_n1079_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X3 a_n487_n500# a_n887_n588# a_n945_n500# a_n1079_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Y9S9FP a_n1174_n500# a_n200_n597# a_200_n500#
+ a_n1116_n597# a_n716_n500# a_n258_n500# w_n1374_n797# a_1116_n500# a_n658_n597#
+ a_658_n500# a_716_n597# a_258_n597#
X0 a_1116_n500# a_716_n597# a_658_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
X1 a_200_n500# a_n200_n597# a_n258_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X2 a_n716_n500# a_n1116_n597# a_n1174_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X3 a_658_n500# a_258_n597# a_200_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X4 a_n258_n500# a_n658_n597# a_n716_n500# w_n1374_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_62W3XE a_358_n500# a_158_n588# a_100_n500# a_n158_n500#
+ a_n358_n588# a_n100_n588# a_n550_n722# a_n416_n500#
X0 a_100_n500# a_n100_n588# a_n158_n500# a_n550_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X1 a_n158_n500# a_n358_n588# a_n416_n500# a_n550_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X2 a_358_n500# a_158_n588# a_100_n500# a_n550_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EC8RE7 a_416_n500# a_n1364_n500# a_830_n588#
+ a_n1676_n722# a_n118_n500# a_1186_n588# a_n594_n588# a_238_n500# a_n1186_n500# a_652_n588#
+ a_1484_n500# a_n830_n500# a_n60_n588# a_950_n500# a_1008_n588# a_n416_n588# a_n1008_n500#
+ a_474_n588# a_n1484_n588# a_n652_n500# a_772_n500# a_n238_n588# a_296_n588# a_n474_n500#
+ a_1128_n500# a_n1306_n588# a_n950_n588# a_594_n500# a_n1542_n500# a_n296_n500# a_118_n588#
+ a_60_n500# a_1364_n588# a_n1128_n588# a_n772_n588#
X0 a_416_n500# a_296_n588# a_238_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 a_n296_n500# a_n416_n588# a_n474_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_1306_n500# a_1186_n588# a_1128_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X3 a_n1364_n500# a_n1484_n588# a_n1542_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X4 a_238_n500# a_118_n588# a_60_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X5 a_1128_n500# a_1008_n588# a_950_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X6 a_n1186_n500# a_n1306_n588# a_n1364_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X7 a_772_n500# a_652_n588# a_594_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_n118_n500# a_n238_n588# a_n296_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X9 a_n652_n500# a_n772_n588# a_n830_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X10 a_n1008_n500# a_n1128_n588# a_n1186_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X11 a_594_n500# a_474_n588# a_416_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X12 a_60_n500# a_n60_n588# a_n118_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X13 a_1484_n500# a_1364_n588# a_1306_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X14 a_950_n500# a_830_n588# a_772_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X15 a_n830_n500# a_n950_n588# a_n1008_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X16 a_n474_n500# a_n594_n588# a_n652_n500# a_n1676_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Y9J9EP a_n358_n597# a_358_n500# a_n100_n597#
+ a_100_n500# a_n158_n500# a_158_n597# w_n616_n797# a_n416_n500#
X0 a_100_n500# a_n100_n597# a_n158_n500# w_n616_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X1 a_n158_n500# a_n358_n597# a_n416_n500# w_n616_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X2 a_358_n500# a_158_n597# a_100_n500# w_n616_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_QZVU2P a_2974_n500# a_2116_n500# a_n458_n500#
+ a_n2974_n588# a_n3032_n500# a_n2116_n588# a_n400_n588# a_1258_n500# a_2174_n588#
+ a_n2174_n500# a_n3166_n722# a_n1258_n588# a_1316_n588# a_458_n588# a_400_n500# a_n1316_n500#
X0 a_n2174_n500# a_n2974_n588# a_n3032_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=4
X1 a_1258_n500# a_458_n588# a_400_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X2 a_n1316_n500# a_n2116_n588# a_n2174_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X3 a_n458_n500# a_n1258_n588# a_n1316_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X4 a_2116_n500# a_1316_n588# a_1258_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X5 a_2974_n500# a_2174_n588# a_2116_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=4
X6 a_400_n500# a_n400_n588# a_n458_n500# a_n3166_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_7JLQGA a_416_n500# a_n238_n597# a_n118_n500#
+ a_296_n597# a_238_n500# a_n830_n500# a_118_n597# a_n772_n597# w_n1030_n797# a_772_n500#
+ a_n474_n500# a_n594_n597# a_652_n597# a_n60_n597# a_n296_n500# a_60_n500# a_n416_n597#
+ a_474_n597#
X0 a_416_n500# a_296_n597# a_238_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X1 a_n296_n500# a_n416_n597# a_n474_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X2 a_238_n500# a_118_n597# a_60_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X3 a_772_n500# a_652_n597# a_594_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.6
X4 a_n118_n500# a_n238_n597# a_n296_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X5 a_n652_n500# a_n772_n597# a_n830_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.6
X6 a_594_n500# a_474_n597# a_416_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X7 a_60_n500# a_n60_n597# a_n118_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
X8 a_n474_n500# a_n594_n597# a_n652_n500# w_n1030_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.6
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_3DCHX4 a_n1687_n1687# a_n3287_n557# a_29_599#
+ a_1629_1781# a_1687_n2869# a_n3287_n1713# a_3287_n2843# a_3287_n531# a_n1629_1755#
+ a_1687_n1713# a_n1687_n531# a_n1687_625# a_29_n2869# a_n3345_n2843# a_n1687_n2843#
+ a_1687_1755# a_29_n1713# a_n29_n531# a_3287_1781# a_29_1755# a_n29_n1687# a_n3345_625#
+ a_n3479_n3003# a_n1687_1781# a_1629_n1687# a_n29_625# a_n3287_1755# a_n1629_n557#
+ a_3287_625# a_1687_599# a_n3345_n531# a_1629_n531# a_n3287_599# a_n1629_n2869# a_3287_n1687#
+ a_n29_1781# a_1629_625# a_n29_n2843# a_1687_n557# a_n1629_n1713# a_n1629_599# a_1629_n2843#
+ a_29_n557# a_n3287_n2869# a_n3345_n1687# a_n3345_1781#
X0 a_1629_1781# a_29_1755# a_n29_1781# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X1 a_3287_n531# a_1687_n557# a_1629_n531# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X2 a_n1687_n531# a_n3287_n557# a_n3345_n531# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X3 a_3287_1781# a_1687_1755# a_1629_1781# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X4 a_n29_625# a_n1629_599# a_n1687_625# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X5 a_n1687_1781# a_n3287_1755# a_n3345_1781# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X6 a_n1687_n1687# a_n3287_n1713# a_n3345_n1687# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X7 a_1629_n1687# a_29_n1713# a_n29_n1687# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X8 a_n1687_n2843# a_n3287_n2869# a_n3345_n2843# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X9 a_3287_n1687# a_1687_n1713# a_1629_n1687# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X10 a_1629_n2843# a_29_n2869# a_n29_n2843# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X11 a_1629_625# a_29_599# a_n29_625# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X12 a_3287_625# a_1687_599# a_1629_625# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X13 a_n29_n531# a_n1629_n557# a_n1687_n531# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X14 a_3287_n2843# a_1687_n2869# a_1629_n2843# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=8
X15 a_n29_1781# a_n1629_1755# a_n1687_1781# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X16 a_n29_n1687# a_n1629_n1713# a_n1687_n1687# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X17 a_n29_n2843# a_n1629_n2869# a_n1687_n2843# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
X18 a_n1687_625# a_n3287_599# a_n3345_625# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=8
X19 a_1629_n531# a_29_n557# a_n29_n531# a_n3479_n3003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_75J6LY a_n3403_n597# a_5977_n500# a_5177_n597#
+ a_29_n597# a_n2603_n500# a_5119_n500# a_n6893_n500# a_3461_n597# a_3403_n500# a_n6035_n500#
+ a_n2545_n597# w_n7093_n797# a_n1745_n500# a_4319_n597# a_n6835_n597# a_2545_n500#
+ a_2603_n597# a_n5177_n500# a_n1687_n597# a_n4261_n597# a_n887_n500# a_6835_n500#
+ a_n3461_n500# a_6035_n597# a_n5977_n597# a_n29_n500# a_n5119_n597# a_1687_n500#
+ a_1745_n597# a_n829_n597# a_4261_n500# a_887_n597# a_829_n500# a_n4319_n500#
X0 a_n29_n500# a_n829_n597# a_n887_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X1 a_n5177_n500# a_n5977_n597# a_n6035_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X2 a_4261_n500# a_3461_n597# a_3403_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X3 a_2545_n500# a_1745_n597# a_1687_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X4 a_n4319_n500# a_n5119_n597# a_n5177_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X5 a_829_n500# a_29_n597# a_n29_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X6 a_n2603_n500# a_n3403_n597# a_n3461_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X7 a_1687_n500# a_887_n597# a_829_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X8 a_6835_n500# a_6035_n597# a_5977_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=4
X9 a_5119_n500# a_4319_n597# a_4261_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X10 a_n3461_n500# a_n4261_n597# a_n4319_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X11 a_n1745_n500# a_n2545_n597# a_n2603_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X12 a_5977_n500# a_5177_n597# a_5119_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X13 a_n887_n500# a_n1687_n597# a_n1745_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
X14 a_n6035_n500# a_n6835_n597# a_n6893_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=4
X15 a_3403_n500# a_2603_n597# a_2545_n500# w_n7093_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=4
.ends

.subckt ibias_gen ibias0 itest ibias1 ibg_200n vbg_1v2 isrc_sel ena ve avss avdd
Xsky130_fd_pr__nfet_g5v0d10v5_XZ4X25_0 isrc_sel_b ena_b isrc_sel avss ena_b vn1 avss
+ avss avss vn0 sky130_fd_pr__nfet_g5v0d10v5_XZ4X25
Xsky130_fd_pr__pfet_g5v0d10v5_Y9S9FP_0 avdd ena vp0 isrc_sel vp1 avdd avdd vp ena
+ avdd ena isrc_sel_b sky130_fd_pr__pfet_g5v0d10v5_Y9S9FP
Xsky130_fd_pr__nfet_g5v0d10v5_62W3XE_0 avss isrc_sel isrc_sel_b ena_b ena avss avss
+ avss sky130_fd_pr__nfet_g5v0d10v5_62W3XE
Xsky130_fd_pr__nfet_g5v0d10v5_EC8RE7_1 vp0 vstart isrc_sel avss vn0 isrc_sel vbg_1v2
+ vn0 vn0 avss ibg_200n vn0 vbg_1v2 vp1 avss vbg_1v2 vstart isrc_sel_b vbg_1v2 vstart
+ vp vbg_1v2 avss vn0 vn1 vbg_1v2 vbg_1v2 vp vn0 vstart vbg_1v2 vstart ena vbg_1v2
+ vbg_1v2 sky130_fd_pr__nfet_g5v0d10v5_EC8RE7
Xsky130_fd_pr__pfet_g5v0d10v5_Y9J9EP_0 ena avdd avdd isrc_sel_b ena_b isrc_sel avdd
+ avdd sky130_fd_pr__pfet_g5v0d10v5_Y9J9EP
Xsky130_fd_pr__nfet_g5v0d10v5_QZVU2P_1 avss vr ve avss avss vn0 avss vp0 avss ve avss
+ vn0 vn0 vn0 vr vn0 sky130_fd_pr__nfet_g5v0d10v5_QZVU2P
Xsky130_fd_pr__res_xhigh_po_1p41_DVQADA_0 m1_4165_119# m1_3409_119# m1_3409_119# m1_5299_7518#
+ m1_1519_7518# m1_385_119# m1_2653_119# m1_385_119# m1_2653_119# m1_6433_119# m1_1897_119#
+ avss m1_6055_7518# m1_3787_7518# m1_2275_7518# m1_1519_7518# m1_6055_7518# m1_4165_119#
+ m1_5299_7518# m1_763_7518# m1_4921_119# m1_763_7518# m1_7189_119# m1_4543_7518#
+ m1_1897_119# m1_7189_119# m1_3031_7518# m1_6811_7518# m1_4921_119# m1_5677_119#
+ m1_5677_119# m1_6811_7518# m1_3031_7518# m1_3787_7518# m1_1141_119# avss m1_4543_7518#
+ m1_1141_119# m1_6433_119# vr m1_2275_7518# sky130_fd_pr__res_xhigh_po_1p41_DVQADA
Xsky130_fd_pr__pfet_g5v0d10v5_7JLQGA_0 vn1 isrc_sel vp avdd vp1 vstart isrc_sel_b
+ ena_b avdd ibg_200n avdd isrc_sel ena_b avdd vp0 vp avdd isrc_sel_b sky130_fd_pr__pfet_g5v0d10v5_7JLQGA
Xsky130_fd_pr__nfet_g5v0d10v5_3DCHX4_0 avss avss vn1 avss avss avss avss avss vn1
+ avss avss avss vn1 avss avss avss vn1 vn1 avss vn1 vp1 avss avss avss avss vp1 avss
+ vn1 avss avss avss avss avss vn1 avss vp1 avss vp1 avss vn1 vn1 avss vn1 avss avss
+ avss sky130_fd_pr__nfet_g5v0d10v5_3DCHX4
Xsky130_fd_pr__pfet_g5v0d10v5_75J6LY_0 vp0 avdd vp vp vp0 ibias1 avdd vp1 vp1 avdd
+ vp0 avdd avdd vp avdd avdd vp1 vn0 avdd avdd avdd avdd avdd avdd vp0 ibias0 vp0
+ itest vp vp avdd vp avdd avdd sky130_fd_pr__pfet_g5v0d10v5_75J6LY
.ends

.subckt sky130_fd_pr__rf_pnp_05v5_W0p68L0p68 Base Collector Emitter m=1
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W0p68L0p68
**devattr s=18496,544
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_T82T27 a_1629_47# a_1687_21# a_n1687_47# a_4945_n309#
+ a_n1629_n335# a_n5137_n469# a_n4945_n335# a_n29_47# a_29_21# a_n3287_21# a_1687_n335#
+ a_3287_n309# a_n5003_n309# a_29_n335# a_n1687_n309# a_n5003_47# a_n4945_21# a_n3287_n335#
+ a_n1629_21# a_3345_21# a_n29_n309# a_3287_47# a_n3345_47# a_3345_n335# a_n3345_n309#
+ a_1629_n309# a_4945_47#
X0 a_n1687_47# a_n3287_21# a_n3345_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1 a_4945_47# a_3345_21# a_3287_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X2 a_1629_n309# a_29_n335# a_n29_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X3 a_n3345_n309# a_n4945_n335# a_n5003_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X4 a_3287_n309# a_1687_n335# a_1629_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X5 a_n1687_n309# a_n3287_n335# a_n3345_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X6 a_n3345_47# a_n4945_21# a_n5003_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X7 a_n29_47# a_n1629_21# a_n1687_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X8 a_4945_n309# a_3345_n335# a_3287_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X9 a_3287_47# a_1687_21# a_1629_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X10 a_n29_n309# a_n1629_n335# a_n1687_n309# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X11 a_1629_47# a_29_21# a_n29_47# a_n5137_n469# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3HV7M9 a_3345_n161# a_n1687_n64# a_n1629_n161#
+ a_n4945_n161# w_n5203_n362# a_1687_n161# a_n3345_n64# a_29_n161# a_3287_n64# a_n29_n64#
+ a_n3287_n161# a_1629_n64# a_n5003_n64# a_4945_n64#
X0 a_n29_n64# a_n1629_n161# a_n1687_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1 a_n3345_n64# a_n4945_n161# a_n5003_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X2 a_1629_n64# a_29_n161# a_n29_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X3 a_3287_n64# a_1687_n161# a_1629_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X4 a_4945_n64# a_3345_n161# a_3287_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X5 a_n1687_n64# a_n3287_n161# a_n3345_n64# w_n5203_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_5H9LZ4 a_n100_n344# a_n158_118# a_n100_21# a_100_n612#
+ a_100_483# a_n100_n709# a_100_n247# a_n158_n612# a_n100_386# a_n158_n247# a_100_118#
+ w_n358_n909# a_n158_483#
X0 a_100_118# a_n100_21# a_n158_118# w_n358_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1 a_100_483# a_n100_386# a_n158_483# w_n358_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 a_100_n612# a_n100_n709# a_n158_n612# w_n358_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_100_n247# a_n100_n344# a_n158_n247# w_n358_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_GG9S2Z a_n100_199# a_100_n487# a_100_581# a_100_n131#
+ a_n158_n487# a_n100_n157# a_n100_555# a_100_n843# a_n158_n131# a_n158_225# a_n100_n869#
+ a_n158_581# a_n158_n843# a_n100_n513# a_n292_n1003# a_100_225#
X0 a_100_n131# a_n100_n157# a_n158_n131# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1 a_100_581# a_n100_555# a_n158_581# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 a_100_n843# a_n100_n869# a_n158_n843# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_100_225# a_n100_199# a_n158_225# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X4 a_100_n487# a_n100_n513# a_n158_n487# a_n292_n1003# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_5HVT2F a_1629_n430# a_4945_n65# a_n3287_n1257#
+ a_n3287_n892# a_3345_n162# a_4945_665# a_n3287_568# w_n5203_n1457# a_3345_n1257#
+ a_3287_1030# a_n1629_933# a_n5003_1030# a_3287_n1160# a_n29_n795# a_n4945_n527#
+ a_n1687_1030# a_3345_933# a_n4945_933# a_1687_n1257# a_4945_n430# a_1687_n527# a_n1629_568#
+ a_29_933# a_29_n527# a_3345_568# a_n4945_568# a_n5003_n1160# a_3345_n892# a_n3345_300#
+ a_n3345_n1160# a_n3345_n795# a_n1687_n65# a_n1629_n162# a_29_568# a_29_n1257# a_1629_n795#
+ a_n3287_n527# a_3287_300# a_n29_300# a_n1687_665# a_n29_1030# a_n1687_n1160# a_3287_n430#
+ a_n5003_n430# a_n1687_n430# a_n4945_n162# a_4945_n795# a_1687_n162# a_1629_300#
+ a_n5003_300# a_n1629_n892# a_1687_203# a_4945_300# a_n3287_203# a_1629_1030# a_n3345_1030#
+ a_3345_n527# a_n3345_n65# a_29_n162# a_n3345_665# a_n4945_n1257# a_n4945_n892# a_n29_n430#
+ a_3287_n65# a_n29_n65# a_n29_665# a_n3287_n162# a_3287_665# a_4945_n1160# a_3287_n795#
+ a_n5003_n795# a_1687_n892# a_n1629_203# a_4945_1030# a_n1629_n1257# a_1687_933#
+ a_n1687_n795# a_3345_203# a_n4945_203# a_n3287_933# a_n29_n1160# a_29_n892# a_1629_n1160#
+ a_n1629_n527# a_1629_n65# a_n5003_n65# a_1629_665# a_n5003_665# a_n3345_n430# a_n1687_300#
+ a_29_203# a_1687_568#
X0 a_n29_300# a_n1629_203# a_n1687_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1 a_3287_n795# a_1687_n892# a_1629_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2 a_n29_1030# a_n1629_933# a_n1687_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X3 a_4945_n430# a_3345_n527# a_3287_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X4 a_n1687_n795# a_n3287_n892# a_n3345_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X5 a_n3345_665# a_n4945_568# a_n5003_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X6 a_n3345_300# a_n4945_203# a_n5003_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X7 a_n1687_n65# a_n3287_n162# a_n3345_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X8 a_n29_n1160# a_n1629_n1257# a_n1687_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X9 a_1629_665# a_29_568# a_n29_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X10 a_4945_n795# a_3345_n892# a_3287_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X11 a_n29_n430# a_n1629_n527# a_n1687_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X12 a_3287_665# a_1687_568# a_1629_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X13 a_1629_1030# a_29_933# a_n29_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X14 a_1629_300# a_29_203# a_n29_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X15 a_4945_665# a_3345_568# a_3287_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X16 a_3287_300# a_1687_203# a_1629_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X17 a_n29_n65# a_n1629_n162# a_n1687_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X18 a_n3345_1030# a_n4945_933# a_n5003_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X19 a_4945_300# a_3345_203# a_3287_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X20 a_3287_1030# a_1687_933# a_1629_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X21 a_n3345_n65# a_n4945_n162# a_n5003_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X22 a_n1687_1030# a_n3287_933# a_n3345_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X23 a_n29_n795# a_n1629_n892# a_n1687_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X24 a_n3345_n1160# a_n4945_n1257# a_n5003_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X25 a_1629_n430# a_29_n527# a_n29_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X26 a_n1687_n1160# a_n3287_n1257# a_n3345_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X27 a_1629_n65# a_29_n162# a_n29_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X28 a_4945_n1160# a_3345_n1257# a_3287_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X29 a_n3345_n430# a_n4945_n527# a_n5003_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X30 a_4945_1030# a_3345_933# a_3287_1030# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X31 a_n1687_665# a_n3287_568# a_n3345_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X32 a_3287_n65# a_1687_n162# a_1629_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X33 a_3287_n430# a_1687_n527# a_1629_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X34 a_1629_n1160# a_29_n1257# a_n29_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X35 a_n1687_300# a_n3287_203# a_n3345_300# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X36 a_4945_n65# a_3345_n162# a_3287_n65# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X37 a_n1687_n430# a_n3287_n527# a_n3345_n430# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X38 a_1629_n795# a_29_n892# a_n29_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X39 a_3287_n1160# a_1687_n1257# a_1629_n1160# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X40 a_n29_665# a_n1629_568# a_n1687_665# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X41 a_n3345_n795# a_n4945_n892# a_n5003_n795# w_n5203_n1457# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_HZHY2Z a_861_n131# a_207_n157# a_n861_n157# a_n563_n131#
+ a_683_n131# a_n919_n131# a_29_n157# a_n683_n157# a_n385_n131# a_n1053_n291# a_741_n157#
+ a_505_n131# a_n505_n157# a_563_n157# a_n207_n131# a_327_n131# a_n327_n157# a_385_n157#
+ a_n29_n131# a_149_n131# a_n741_n131# a_n149_n157#
X0 a_505_n131# a_385_n157# a_327_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X1 a_n385_n131# a_n505_n157# a_n563_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2 a_327_n131# a_207_n157# a_149_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X3 a_149_n131# a_29_n157# a_n29_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X4 a_861_n131# a_741_n157# a_683_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X5 a_n207_n131# a_n327_n157# a_n385_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X6 a_n741_n131# a_n861_n157# a_n919_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X7 a_683_n131# a_563_n157# a_505_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X8 a_n29_n131# a_n149_n157# a_n207_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X9 a_n563_n131# a_n683_n157# a_n741_n131# a_n1053_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ZV8547 a_3345_439# a_3287_527# a_1687_21# a_n4945_439#
+ a_n5003_n1563# a_1629_n1145# a_3345_n815# a_3287_n727# a_29_439# a_n5003_n727# a_n3345_n1563#
+ a_n4945_1275# a_n29_1363# a_4945_n309# a_3345_n397# a_n1687_n727# a_1687_1275# a_n1687_n1563#
+ a_n5003_527# a_1629_527# a_n4945_n1651# a_29_n1233# a_3287_n1145# a_n3345_109# a_29_1275#
+ a_4945_527# a_n1687_945# a_n3287_21# a_n29_109# a_3287_109# a_n3345_1363# a_29_21#
+ a_n5003_n1145# a_n1629_n1651# a_n1629_n815# a_1629_1363# a_n3287_1275# a_1687_857#
+ a_3287_n309# a_n29_n727# a_n5003_n309# a_n3345_n1145# a_n3287_857# a_n1629_n397#
+ a_n1687_n309# a_n1687_n1145# a_n5003_109# a_1629_109# a_n4945_n815# a_n4945_n1233#
+ a_n3287_n1651# a_4945_1363# a_n4945_21# a_4945_n1563# a_n3345_945# a_1687_n815#
+ a_3345_n1651# a_n1629_21# a_4945_109# a_n1687_527# a_n4945_n397# a_n3345_n727# a_n1629_857#
+ a_3345_1275# a_n29_n1563# a_1629_n727# a_1687_n1651# a_29_n815# a_n29_945# a_n1629_n1233#
+ a_1687_n397# a_3345_857# a_3287_945# a_n4945_857# a_3345_21# a_1629_n1563# a_1687_439#
+ a_n29_n309# a_29_n397# a_29_857# a_n3287_439# a_n3287_n815# a_3287_1363# a_n5003_1363#
+ a_4945_n727# a_n5137_n1785# a_n3287_n1233# a_n1687_1363# a_n5003_945# a_1629_945#
+ a_4945_n1145# a_29_n1651# a_3287_n1563# a_n3345_527# a_n3287_n397# a_3345_n1233#
+ a_4945_945# a_n1687_109# a_n1629_1275# a_n3345_n309# a_n1629_439# a_n29_n1145# a_1629_n309#
+ a_1687_n1233# a_n29_527#
X0 a_3287_945# a_1687_857# a_1629_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X1 a_1629_109# a_29_21# a_n29_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X2 a_3287_109# a_1687_21# a_1629_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X3 a_4945_n727# a_3345_n815# a_3287_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X4 a_4945_945# a_3345_857# a_3287_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X5 a_4945_109# a_3345_21# a_3287_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X6 a_n29_527# a_n1629_439# a_n1687_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X7 a_n29_1363# a_n1629_1275# a_n1687_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X8 a_n3345_n1145# a_n4945_n1233# a_n5003_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X9 a_1629_n309# a_29_n397# a_n29_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X10 a_n1687_n1145# a_n3287_n1233# a_n3345_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X11 a_n3345_527# a_n4945_439# a_n5003_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X12 a_4945_n1145# a_3345_n1233# a_3287_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X13 a_n29_n1563# a_n1629_n1651# a_n1687_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X14 a_n3345_n309# a_n4945_n397# a_n5003_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X15 a_3287_n309# a_1687_n397# a_1629_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X16 a_n29_n727# a_n1629_n815# a_n1687_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X17 a_1629_n1145# a_29_n1233# a_n29_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X18 a_n1687_n309# a_n3287_n397# a_n3345_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X19 a_n1687_945# a_n3287_857# a_n3345_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X20 a_1629_527# a_29_439# a_n29_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X21 a_n1687_109# a_n3287_21# a_n3345_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X22 a_3287_n1145# a_1687_n1233# a_1629_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X23 a_1629_1363# a_29_1275# a_n29_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X24 a_3287_527# a_1687_439# a_1629_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X25 a_4945_527# a_3345_439# a_3287_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X26 a_4945_n309# a_3345_n397# a_3287_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X27 a_n3345_1363# a_n4945_1275# a_n5003_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X28 a_n29_945# a_n1629_857# a_n1687_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X29 a_3287_1363# a_1687_1275# a_1629_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X30 a_n3345_n1563# a_n4945_n1651# a_n5003_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X31 a_n29_109# a_n1629_21# a_n1687_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X32 a_1629_n727# a_29_n815# a_n29_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X33 a_n1687_1363# a_n3287_1275# a_n3345_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X34 a_n1687_n1563# a_n3287_n1651# a_n3345_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X35 a_4945_n1563# a_3345_n1651# a_3287_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X36 a_n3345_945# a_n4945_857# a_n5003_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X37 a_n3345_n727# a_n4945_n815# a_n5003_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X38 a_n3345_109# a_n4945_21# a_n5003_109# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X39 a_3287_n727# a_1687_n815# a_1629_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X40 a_n29_n1145# a_n1629_n1233# a_n1687_n1145# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X41 a_n1687_n727# a_n3287_n815# a_n3345_n727# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X42 a_1629_n1563# a_29_n1651# a_n29_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X43 a_n29_n309# a_n1629_n397# a_n1687_n309# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X44 a_4945_1363# a_3345_1275# a_3287_1363# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X45 a_1629_945# a_29_857# a_n29_945# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X46 a_n1687_527# a_n3287_439# a_n3345_527# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X47 a_3287_n1563# a_1687_n1651# a_1629_n1563# a_n5137_n1785# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_5HV9F5 a_1629_118# a_n5003_118# a_1687_21# a_n29_n612#
+ a_n3287_n344# a_4945_118# a_29_386# a_n1687_483# a_n29_n247# a_n3345_n612# a_n1629_n709#
+ a_1629_n612# a_3345_n344# a_29_21# a_n3287_21# a_n3345_n247# a_n3345_483# w_n5203_n909#
+ a_n4945_n709# a_1629_n247# a_4945_n612# a_n1687_118# a_1687_n709# a_3287_483# a_n29_483#
+ a_29_n709# a_n4945_21# a_n1629_21# a_4945_n247# a_n1629_n344# a_n3287_n709# a_1629_483#
+ a_n5003_483# a_3345_21# a_1687_386# a_3287_n612# a_n5003_n612# a_n3345_118# a_4945_483#
+ a_n3287_386# a_n1687_n612# a_n4945_n344# a_n29_118# a_3287_n247# a_n5003_n247# a_1687_n344#
+ a_3287_118# a_n1687_n247# a_n1629_386# a_3345_n709# a_29_n344# a_3345_386# a_n4945_386#
X0 a_4945_n247# a_3345_n344# a_3287_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X1 a_4945_n612# a_3345_n709# a_3287_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X2 a_n29_118# a_n1629_21# a_n1687_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X3 a_n1687_483# a_n3287_386# a_n3345_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X4 a_n3345_118# a_n4945_21# a_n5003_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X5 a_n29_483# a_n1629_386# a_n1687_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X6 a_n29_n247# a_n1629_n344# a_n1687_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X7 a_n29_n612# a_n1629_n709# a_n1687_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X8 a_1629_118# a_29_21# a_n29_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X9 a_n3345_483# a_n4945_386# a_n5003_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X10 a_3287_118# a_1687_21# a_1629_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X11 a_4945_118# a_3345_21# a_3287_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X12 a_1629_483# a_29_386# a_n29_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X13 a_1629_n612# a_29_n709# a_n29_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X14 a_3287_483# a_1687_386# a_1629_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X15 a_1629_n247# a_29_n344# a_n29_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X16 a_n3345_n247# a_n4945_n344# a_n5003_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X17 a_n3345_n612# a_n4945_n709# a_n5003_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=8
X18 a_4945_483# a_3345_386# a_3287_483# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=8
X19 a_3287_n247# a_1687_n344# a_1629_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X20 a_3287_n612# a_1687_n709# a_1629_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X21 a_n1687_n247# a_n3287_n344# a_n3345_n247# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X22 a_n1687_n612# a_n3287_n709# a_n3345_n612# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
X23 a_n1687_118# a_n3287_21# a_n3345_118# w_n5203_n909# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_W8MWAU a_n741_n136# w_n1119_n362# a_861_n136#
+ a_n327_n162# a_385_n162# a_n563_n136# a_683_n136# a_n149_n162# a_n919_n136# a_207_n162#
+ a_n385_n136# a_n861_n162# a_505_n136# a_29_n162# a_n207_n136# a_n683_n162# a_741_n162#
+ a_327_n136# a_n505_n162# a_n29_n136# a_563_n162# a_149_n136#
X0 a_861_n136# a_741_n162# a_683_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.6
X1 a_n207_n136# a_n327_n162# a_n385_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X2 a_n741_n136# a_n861_n162# a_n919_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.6
X3 a_683_n136# a_563_n162# a_505_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X4 a_n29_n136# a_n149_n162# a_n207_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X5 a_n563_n136# a_n683_n162# a_n741_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X6 a_505_n136# a_385_n162# a_327_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X7 a_n385_n136# a_n505_n162# a_n563_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X8 a_327_n136# a_207_n162# a_149_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
X9 a_149_n136# a_29_n162# a_n29_n136# w_n1119_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.6
.ends

.subckt comparator ibias out ena vinn vinp avss vt avdd
Xsky130_fd_pr__nfet_g5v0d10v5_T82T27_1 n0 vm vm avss vn avss avss avss vm vm vn avss
+ avss vn vn avss avss vn vm avss avss avss avss avss avss vt avss sky130_fd_pr__nfet_g5v0d10v5_T82T27
Xsky130_fd_pr__pfet_g5v0d10v5_3HV7M9_0 avdd vm vnn avdd avdd vpp avdd vpp avdd avdd
+ vnn n0 avdd avdd sky130_fd_pr__pfet_g5v0d10v5_3HV7M9
Xsky130_fd_pr__pfet_g5v0d10v5_5H9LZ4_0 ena avdd ena vn vpp ena_b ena_b ibias ena avdd
+ vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5_5H9LZ4
Xsky130_fd_pr__nfet_g5v0d10v5_GG9S2Z_0 ena vm vn vn avss ena_b ena n0 avss avss ena_b
+ ibias avss ena_b avss ena_b sky130_fd_pr__nfet_g5v0d10v5_GG9S2Z
Xsky130_fd_pr__pfet_g5v0d10v5_5HVT2F_0 vnn avdd vnn vnn avdd avdd vnn avdd avdd avdd
+ vnn avdd avdd avdd avdd vpp avdd avdd vpp avdd vpp vnn vpp vpp avdd avdd avdd avdd
+ avdd avdd avdd vpp vnn vpp vpp vnn vnn avdd avdd vpp avdd vpp avdd avdd vpp avdd
+ avdd vpp vnn avdd vnn vpp avdd vnn vnn avdd avdd avdd vpp avdd avdd avdd avdd avdd
+ avdd avdd vnn avdd avdd avdd avdd vpp vnn avdd vnn vpp vpp avdd avdd vnn avdd vpp
+ vnn vnn vnn avdd vnn avdd avdd vpp vpp vpp sky130_fd_pr__pfet_g5v0d10v5_5HVT2F
Xsky130_fd_pr__nfet_g5v0d10v5_HZHY2Z_0 avss n1 n1 avss n1 avss n1 n1 out avss n0 avss
+ n1 n0 avss out n1 n1 out avss out n1 sky130_fd_pr__nfet_g5v0d10v5_HZHY2Z
Xsky130_fd_pr__nfet_g5v0d10v5_ZV8547_0 avss vnn vinn avss vt vt avss vnn vinp vt vnn
+ avss vpp vt avss vt vinn vt vt vt avss vinp vnn vnn vinp vt vt vinn vpp vnn vnn
+ vinp vt vinp vinp vt vinn vinn vnn vpp vt vnn vinn vinp vt vt vt vt avss avss vinn
+ vt avss vt vnn vinn avss vinp vt vt avss vnn vinp avss vpp vt vinn vinp vpp vinp
+ vinn avss vnn avss avss vt vinn vpp vinp vinp vinn vinn vnn vt vt vt vinn vt vt
+ vt vt vinp vnn vnn vinn avss vt vt vinp vnn vinp vpp vt vinn vpp sky130_fd_pr__nfet_g5v0d10v5_ZV8547
Xsky130_fd_pr__pfet_g5v0d10v5_5HV9F5_0 vnn avdd vnn avdd vpp avdd vnn vpp avdd avdd
+ vpp vnn avdd vnn vpp avdd avdd avdd avdd vnn avdd vpp vnn avdd avdd vnn avdd vpp
+ avdd vpp vpp vnn avdd avdd vnn avdd avdd avdd avdd vpp vpp avdd avdd avdd avdd vnn
+ avdd vpp vpp avdd vnn avdd avdd sky130_fd_pr__pfet_g5v0d10v5_5HV9F5
Xsky130_fd_pr__pfet_g5v0d10v5_W8MWAU_0 out avdd avdd n1 n1 avdd n1 n1 avdd n1 out
+ n1 avdd n1 avdd n1 n0 out n1 out n0 avdd sky130_fd_pr__pfet_g5v0d10v5_W8MWAU
.ends

.subckt brownout_ana otrip_decoded[7] otrip_decoded[5] otrip_decoded[3] otrip_decoded[1]
+ vin_vunder vbg_1v2 ena ibg_200n itest isrc_sel vtrip_decoded[7] vtrip_decoded[6]
+ vtrip_decoded[5] vtrip_decoded[4] vtrip_decoded[3] vtrip_decoded[2] vtrip_decoded[0]
+ dcomp brout_filt osc_ena vunder outb comparator_1/vt otrip_decoded[4] dvdd comparator_0/vt
+ otrip_decoded[2] osc_ck outb_unbuf avdd vtrip_decoded[1] otrip_decoded[6] otrip_decoded[0]
+ vin_brout avss dvss
Xsky130_fd_sc_hd__inv_16_3 sky130_fd_sc_hd__inv_4_4/Y dvss dvss dvdd dvdd outb sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hvl__lsbufhv2lv_1_0 dcomp3v3 dvdd dvss avdd avdd vl avdd dvss dvss sky130_fd_sc_hvl__lsbufhv2lv_1
Xsky130_fd_sc_hvl__lsbufhv2lv_1_1 dcomp3v3uv dvdd dvss avdd avdd sky130_fd_sc_hd__inv_4_2/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbufhv2lv_1
Xrstring_mux_0 vin_brout ibias_gen_0/ena rstring_mux_0/otrip_decoded_avdd[7] rstring_mux_0/otrip_decoded_avdd[6]
+ rstring_mux_0/otrip_decoded_avdd[5] rstring_mux_0/otrip_decoded_avdd[4] rstring_mux_0/otrip_decoded_avdd[3]
+ rstring_mux_0/otrip_decoded_avdd[2] rstring_mux_0/otrip_decoded_avdd[1] rstring_mux_0/vtrip_decoded_avdd[7]
+ rstring_mux_0/vtrip_decoded_avdd[6] rstring_mux_0/vtrip_decoded_avdd[5] rstring_mux_0/vtrip_decoded_avdd[4]
+ rstring_mux_0/vtrip_decoded_avdd[3] rstring_mux_0/vtrip_decoded_avdd[2] rstring_mux_0/vtrip_decoded_avdd[1]
+ rstring_mux_0/vtrip_decoded_avdd[0] vin_vunder rstring_mux_0/vtop rstring_mux_0/otrip_decoded_avdd[0]
+ avdd avss rstring_mux
Xsky130_fd_sc_hd__inv_4_0 schmitt_trigger_0/out dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_0/Y
+ sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_4_1 sky130_fd_sc_hd__inv_4_2/Y dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_1/Y
+ sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_4_2 sky130_fd_sc_hd__inv_4_2/A dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_2/Y
+ sky130_fd_sc_hd__inv_4
Xschmitt_trigger_0 schmitt_trigger_0/in schmitt_trigger_0/out dvdd dvss schmitt_trigger
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|0] otrip_decoded[0] dvdd dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[0]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|0] otrip_decoded[1] dvdd dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[1]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|1] otrip_decoded[2] dvdd dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[2]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|1] otrip_decoded[3] dvdd dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[3]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|2] otrip_decoded[4] dvdd dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[4]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|2] otrip_decoded[5] dvdd dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[5]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|3] otrip_decoded[6] dvdd dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[6]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|3] otrip_decoded[7] dvdd dvss avdd avdd rstring_mux_0/otrip_decoded_avdd[7]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|4] vtrip_decoded[0] dvdd dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[0]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|4] vtrip_decoded[1] dvdd dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[1]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|5] vtrip_decoded[2] dvdd dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[2]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|5] vtrip_decoded[3] dvdd dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[3]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|6] vtrip_decoded[4] dvdd dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[4]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6] vtrip_decoded[5] dvdd dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[5]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|7] vtrip_decoded[6] dvdd dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[6]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|7] vtrip_decoded[7] dvdd dvss avdd avdd rstring_mux_0/vtrip_decoded_avdd[7]
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|8] ena dvdd dvss avdd avdd ibias_gen_0/ena avdd
+ dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|8] isrc_sel dvdd dvss avdd avdd ibias_gen_0/isrc_sel
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xrc_osc_0 dvdd osc_ck osc_ena dvss rc_osc
Xsky130_fd_sc_hd__inv_4_3 vl dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_3/Y sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_4_4 outb_unbuf dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_4_4/Y
+ sky130_fd_sc_hd__inv_4
Xsky130_fd_pr__res_xhigh_po_1p41_DVQADA_0 m1_n11325_2001# m1_n11325_2001# m1_n12081_2001#
+ m1_n10191_9400# m1_n13971_9400# m1_n14349_2001# m1_n12081_2001# vl m1_n12837_2001#
+ m1_n8301_2001# m1_n12837_2001# avss m1_n9435_9400# m1_n10947_9400# m1_n13215_9400#
+ m1_n13215_9400# m1_n8679_9400# m1_n10569_2001# m1_n9435_9400# m1_n13971_9400# m1_n10569_2001#
+ m1_n14727_9400# m1_n8301_2001# m1_n10947_9400# m1_n13593_2001# schmitt_trigger_0/in
+ m1_n11703_9400# m1_n8679_9400# m1_n9813_2001# m1_n9057_2001# m1_n9813_2001# m1_n7923_9400#
+ m1_n12459_9400# m1_n11703_9400# m1_n13593_2001# m1_n14727_9400# m1_n10191_9400#
+ m1_n14349_2001# m1_n9057_2001# m1_n7923_9400# m1_n12459_9400# sky130_fd_pr__res_xhigh_po_1p41_DVQADA
Xsky130_fd_pr__cap_mim_m3_2_LUWKLG_0 schmitt_trigger_0/in dvss sky130_fd_pr__cap_mim_m3_2_LUWKLG
Xibias_gen_0 ibias_gen_0/ibias0 itest ibias_gen_0/ibias1 ibg_200n vbg_1v2 ibias_gen_0/isrc_sel
+ ibias_gen_0/ena ibias_gen_0/ve avss avdd ibias_gen
Xsky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0 avss avss ibias_gen_0/ve sky130_fd_pr__rf_pnp_05v5_W0p68L0p68 m=1
Xcomparator_0 ibias_gen_0/ibias1 dcomp3v3uv ibias_gen_0/ena vin_vunder vbg_1v2 avss
+ comparator_0/vt avdd comparator
Xcomparator_1 ibias_gen_0/ibias0 dcomp3v3 ibias_gen_0/ena vin_brout vbg_1v2 avss comparator_1/vt
+ avdd comparator
Xsky130_fd_sc_hd__inv_16_0 sky130_fd_sc_hd__inv_4_0/Y dvss dvss dvdd dvdd brout_filt
+ sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_1 sky130_fd_sc_hd__inv_4_1/Y dvss dvss dvdd dvdd vunder sky130_fd_sc_hd__inv_16
Xsky130_fd_sc_hd__inv_16_2 sky130_fd_sc_hd__inv_4_3/Y dvss dvss dvdd dvdd dcomp sky130_fd_sc_hd__inv_16
.ends

.subckt sky130_ajc_ip__brownout avdd outb dvdd osc_ck dcomp vbg_1v2 otrip[2] otrip[1]
+ otrip[0] itest brout_filt vtrip[2] vtrip[1] vtrip[0] vin_brout ena force_ena_rc_osc
+ vin_vunder force_dis_rc_osc timed_out vunder force_short_oneshot isrc_sel ibg_200n
+ brownout_ana_0/comparator_1/vt brownout_ana_0/comparator_0/vt avss dvss
Xsky130_fd_pr__nfet_g5v0d10v5_PXF6AN_0 dvss dvss ena dvss dvss dvss dvss dvss dvss
+ dvss otrip[1] dvss dvss force_short_oneshot dvss dvss dvss dvss dvss force_dis_rc_osc
+ dvss otrip[2] force_ena_rc_osc dvss dvss dvss dvss otrip[0] isrc_sel dvss dvss dvss
+ dvss dvss sky130_fd_pr__nfet_g5v0d10v5_PXF6AN
Xbrownout_dig_0 dvdd brout_filt dcomp ena force_dis_rc_osc force_ena_rc_osc force_short_oneshot
+ osc_ck otrip[0] otrip[1] otrip[2] vtrip[0] vtrip[1] vtrip[2] brownout_dig_0/osc_ena
+ brownout_dig_0/otrip_decoded[0] brownout_dig_0/otrip_decoded[1] brownout_dig_0/otrip_decoded[3]
+ brownout_dig_0/otrip_decoded[4] brownout_dig_0/otrip_decoded[5] brownout_dig_0/otrip_decoded[6]
+ brownout_dig_0/otrip_decoded[7] brownout_dig_0/outb_unbuf timed_out brownout_dig_0/vtrip_decoded[0]
+ brownout_dig_0/vtrip_decoded[1] brownout_dig_0/vtrip_decoded[2] brownout_dig_0/vtrip_decoded[3]
+ brownout_dig_0/vtrip_decoded[4] brownout_dig_0/vtrip_decoded[5] brownout_dig_0/vtrip_decoded[6]
+ brownout_dig_0/vtrip_decoded[7] brownout_dig_0/otrip_decoded[2] dvss brownout_dig
Xsky130_fd_pr__nfet_g5v0d10v5_V6EN4F_0 dvss vin_vunder dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_V6EN4F
Xsky130_fd_pr__nfet_g5v0d10v5_XTZQRT_0 dvss dvss vtrip[1] dvss dvss dvss dvss dvss
+ dvss dvss vin_brout dvss dvss dvss dvss vbg_1v2 vtrip[2] dvss dvss dvss vtrip[0]
+ dvss sky130_fd_pr__nfet_g5v0d10v5_XTZQRT
Xbrownout_ana_0 brownout_dig_0/otrip_decoded[7] brownout_dig_0/otrip_decoded[5] brownout_dig_0/otrip_decoded[3]
+ brownout_dig_0/otrip_decoded[1] vin_vunder vbg_1v2 ena ibg_200n itest isrc_sel brownout_dig_0/vtrip_decoded[7]
+ brownout_dig_0/vtrip_decoded[6] brownout_dig_0/vtrip_decoded[5] brownout_dig_0/vtrip_decoded[4]
+ brownout_dig_0/vtrip_decoded[3] brownout_dig_0/vtrip_decoded[2] brownout_dig_0/vtrip_decoded[0]
+ dcomp brout_filt brownout_dig_0/osc_ena vunder outb brownout_ana_0/comparator_1/vt
+ brownout_dig_0/otrip_decoded[4] dvdd brownout_ana_0/comparator_0/vt brownout_dig_0/otrip_decoded[2]
+ osc_ck brownout_dig_0/outb_unbuf avdd brownout_dig_0/vtrip_decoded[1] brownout_dig_0/otrip_decoded[6]
+ brownout_dig_0/otrip_decoded[0] vin_brout avss dvss brownout_ana
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_BWAZV5 a_n700_n197# a_700_n100# w_n958_n397#
+ a_n758_n100#
X0 a_700_n100# a_n700_n197# a_n758_n100# w_n958_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=7
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_A2FZRM a_n900_n188# a_n900_n1024# a_900_n518#
+ a_n900_648# a_n958_318# a_n958_n518# a_900_736# a_n1102_n1158# a_900_n100# a_900_n936#
+ a_900_318# a_n900_230# a_n958_n100# a_n958_736# a_n958_n936# a_n900_n606#
X0 a_900_n100# a_n900_n188# a_n958_n100# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
X1 a_900_n518# a_n900_n606# a_n958_n518# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
X2 a_900_318# a_n900_230# a_n958_318# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
X3 a_900_n936# a_n900_n1024# a_n958_n936# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
X4 a_900_736# a_n900_648# a_n958_736# a_n1102_n1158# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=9
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0 a_n252_n322# a_50_n100# a_n108_n100#
+ a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n252_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLAZY6__0 a_n50_n197# a_50_n100# w_n308_n397#
+ a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n308_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_PC2PN5 w_n1258_n397# a_n1000_n197# a_1000_n100#
+ a_n1058_n100#
X0 a_1000_n100# a_n1000_n197# a_n1058_n100# w_n1258_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_69K6TN a_700_n100# a_n758_n100# a_n700_n188#
+ a_n902_n322#
X0 a_700_n100# a_n700_n188# a_n758_n100# a_n902_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=7
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_QZEXQH a_1044_n1416# a_214_n1416# a_n1114_n1416#
+ a_546_984# a_n1114_984# a_n118_984# a_48_n1416# a_1376_n1416# a_n450_984# a_n782_n1416#
+ a_878_984# a_546_n1416# a_n1446_984# a_712_984# a_n1446_n1416# a_n284_n1416# a_n616_n1416#
+ a_n782_984# a_1210_n1416# a_1044_984# a_878_n1416# a_n118_n1416# a_n616_984# a_48_984#
+ a_380_984# a_1376_984# a_n948_n1416# a_n1576_n1546# a_380_n1416# a_n948_984# a_712_n1416#
+ a_1210_984# a_214_984# a_n1280_n1416# a_n284_984# a_n450_n1416# a_n1280_984#
X0 a_n118_984# a_n118_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X1 a_n1280_984# a_n1280_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X2 a_n948_984# a_n948_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X3 a_1210_984# a_1210_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X4 a_n616_984# a_n616_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X5 a_380_984# a_380_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X6 a_878_984# a_878_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X7 a_546_984# a_546_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X8 a_n1446_984# a_n1446_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X9 a_214_984# a_214_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X10 a_1376_984# a_1376_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X11 a_n1114_984# a_n1114_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X12 a_n284_984# a_n284_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X13 a_1044_984# a_1044_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X14 a_n450_984# a_n450_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X15 a_48_984# a_48_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X16 a_712_984# a_712_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X17 a_n782_984# a_n782_n1416# a_n1576_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_Z7JM9H a_1044_n1416# a_214_n1416# a_n2276_984#
+ a_n2110_n1416# a_1542_984# a_n1114_n1416# a_2870_n1416# a_546_984# a_n1114_984#
+ a_n118_984# a_n2110_984# a_1874_n1416# a_2538_984# a_48_n1416# a_n2940_n1416# a_2372_n1416#
+ a_n1944_n1416# a_1874_984# a_n782_n1416# a_n450_984# a_1376_n1416# a_2870_984# a_878_984#
+ a_2704_n1416# a_546_n1416# a_n1446_984# a_n2442_984# a_1708_n1416# a_n2442_n1416#
+ a_n1446_n1416# a_712_984# a_n284_n1416# a_1708_984# a_2206_n1416# a_2704_984# a_n782_984#
+ a_n616_n1416# a_n1778_984# a_n2774_984# a_1210_n1416# a_1044_984# a_2040_984# a_n1612_984#
+ a_878_n1416# a_n118_n1416# a_n616_984# a_n2774_n1416# a_n2608_984# a_n1778_n1416#
+ a_48_984# a_2538_n1416# a_380_984# a_1376_984# a_n948_n1416# a_2372_984# a_n1944_984#
+ a_380_n1416# a_n2276_n1416# a_n948_984# a_n3070_n1546# a_n2940_984# a_1542_n1416#
+ a_712_n1416# a_n2608_n1416# a_1210_984# a_n1280_n1416# a_214_984# a_2040_n1416#
+ a_n1612_n1416# a_n1280_984# a_2206_984# a_n450_n1416# a_n284_984#
X0 a_n2276_984# a_n2276_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X1 a_n118_984# a_n118_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X2 a_1542_984# a_1542_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X3 a_n1280_984# a_n1280_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X4 a_n948_984# a_n948_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X5 a_2704_984# a_2704_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X6 a_1210_984# a_1210_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X7 a_1708_984# a_1708_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X8 a_n616_984# a_n616_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X9 a_380_984# a_380_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X10 a_n2774_984# a_n2774_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X11 a_n2110_984# a_n2110_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X12 a_878_984# a_878_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X13 a_n1778_984# a_n1778_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X14 a_n2442_984# a_n2442_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X15 a_n2940_984# a_n2940_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X16 a_546_984# a_546_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X17 a_n1446_984# a_n1446_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X18 a_2372_984# a_2372_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X19 a_214_984# a_214_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X20 a_1376_984# a_1376_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X21 a_n2608_984# a_n2608_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X22 a_n1114_984# a_n1114_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X23 a_n284_984# a_n284_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X24 a_2040_984# a_2040_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X25 a_2538_984# a_2538_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X26 a_1044_984# a_1044_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X27 a_n1944_984# a_n1944_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X28 a_n450_984# a_n450_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X29 a_48_984# a_48_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X30 a_2206_984# a_2206_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X31 a_2870_984# a_2870_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X32 a_712_984# a_712_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X33 a_1874_984# a_1874_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X34 a_n1612_984# a_n1612_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
X35 a_n782_984# a_n782_n1416# a_n3070_n1546# sky130_fd_pr__res_xhigh_po_0p35 l=10
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_743D3R a_n248_n2546# a_48_n2416# a_n118_1984#
+ a_n118_n2416# a_48_1984#
X0 a_48_1984# a_48_n2416# a_n248_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
X1 a_n118_1984# a_n118_n2416# a_n248_n2546# sky130_fd_pr__res_xhigh_po_0p35 l=20
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MRZGNS c1_n1646_n1500# m3_n1686_n1540#
X0 c1_n1646_n1500# m3_n1686_n1540# sky130_fd_pr__cap_mim_m3_1 l=15 w=15
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_VCAG9S__0 m3_n686_n540# c1_n646_n500#
X0 c1_n646_n500# m3_n686_n540# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PXBJUB a_n1000_n188# a_n1192_n322# a_1000_n100#
+ a_n1058_n100#
X0 a_1000_n100# a_n1000_n188# a_n1058_n100# a_n1192_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_47NWVV a_n258_n100# a_n200_n197# a_200_n100#
+ w_n458_n397#
X0 a_200_n100# a_n200_n197# a_n258_n100# w_n458_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=2
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_YHRXVR a_n129_n2415# a_819_2457# a_n977_2545#
+ a_n1609_n4763# a_n1135_n1109# a_n1551_21# a_n503_n4763# a_603_n3545# a_1235_109#
+ a_n1609_n1109# a_n29_4981# a_445_3763# a_n1135_109# a_n1077_2457# a_n1235_n2415#
+ a_n503_n1109# a_1393_4981# a_n29_1327# a_345_2457# a_1235_n3545# a_977_n3633# a_n761_3675#
+ a_n603_n2415# a_1393_1327# a_1293_3675# a_n919_2457# a_977_21# a_n345_n4763# a_445_n3545#
+ a_n503_2545# a_129_2545# a_n1077_n2415# a_n187_4981# a_n1293_2545# a_n819_n4763#
+ a_919_n3545# a_n345_n1109# a_n1551_3675# a_187_21# a_1077_3763# a_n1451_n4763# a_29_n4851#
+ a_1077_n3545# a_977_2457# a_n187_1327# a_n819_n1109# a_503_n2415# a_n129_n1197#
+ a_n445_n2415# a_n445_2457# a_n1451_n1109# a_n977_109# a_1077_109# a_n919_n2415#
+ a_n1235_n1197# a_1135_n2415# a_n1551_n2415# a_29_4893# a_n187_n4763# a_287_n3545#
+ a_1451_21# a_29_1239# a_1551_n3545# a_n187_n1109# a_603_3763# a_n603_n1197# a_n1293_n4763#
+ a_n1235_2457# a_n129_4893# a_345_n2415# a_1551_4981# a_n287_n2415# a_129_109# a_n1293_n1109#
+ a_n129_1239# a_503_2457# a_n661_2545# a_n445_21# a_819_n2415# a_29_n6069# a_287_2545#
+ a_n661_n4763# a_761_n3545# a_1551_1327# a_n819_4981# a_n29_n3545# a_187_4893# a_1451_3675#
+ a_n1077_n1197# a_n1393_n2415# a_n661_n1109# a_n819_1327# a_187_1239# a_1393_n3545#
+ a_503_n1197# a_n445_n1197# a_n761_n2415# a_n345_4981# a_n1451_2545# a_187_n2415#
+ a_n919_n1197# a_n1609_109# a_n1609_4981# a_1235_3763# a_1135_n1197# a_n345_1327#
+ a_n1551_n1197# a_1451_n2415# a_n603_2457# a_n1609_1327# a_129_n5981# a_1135_2457#
+ a_n1077_21# a_761_3763# a_n977_n4763# a_n1393_2457# a_n287_4893# a_129_n2327# a_345_n1197#
+ a_n1135_4981# a_n977_n1109# a_661_n2415# a_n287_1239# a_661_2457# a_n29_109# a_n287_n1197#
+ a_919_2545# a_1551_109# a_819_n1197# a_n129_n4851# a_819_4893# a_n1135_1327# a_n977_4981#
+ a_n1451_109# a_n1135_n3545# a_345_21# a_29_21# a_n1393_n1197# a_1293_n2415# a_603_n5981#
+ a_819_1239# a_n977_1327# a_n1609_n3545# a_n1077_4893# a_n1235_n4851# a_603_n2327#
+ a_n503_n3545# a_n29_3763# a_445_2545# a_n1077_1239# a_n503_109# a_n761_n1197# a_1235_n5981#
+ a_345_4893# a_187_n1197# a_1393_3763# a_n603_n4851# a_603_109# a_345_1239# a_1235_n2327#
+ a_1451_n1197# a_977_n2415# a_n761_2457# a_1293_2457# a_n919_4893# a_n503_4981# a_445_n5981#
+ a_129_4981# a_n1077_n4851# a_n129_n6069# a_n1293_4981# a_n919_1239# a_919_n5981#
+ a_n503_1327# a_n603_21# a_445_n2327# a_n345_n3545# a_661_n1197# a_129_1327# a_1077_n5981#
+ a_n187_3763# a_n1293_1327# a_1393_109# a_n819_n3545# a_977_4893# a_919_n2327# a_503_n4851#
+ a_n1293_109# a_n1235_n6069# a_n445_n4851# a_n1551_2457# a_1077_2545# a_n445_4893#
+ a_29_n3633# a_n1451_n3545# a_1077_n2327# a_977_1239# a_1293_n1197# a_n919_n4851#
+ a_n445_1239# a_1135_n4851# a_n1551_n4851# a_n603_n6069# a_287_n5981# a_n345_109#
+ a_29_3675# a_1551_n5981# a_287_n2327# a_n187_n3545# a_445_109# a_n1235_4893# a_1551_n2327#
+ a_345_n4851# a_977_n1197# a_n1077_n6069# a_n287_n4851# a_n1235_21# a_603_2545# a_n129_3675#
+ a_n1235_1239# a_n1293_n3545# a_503_4893# a_n661_4981# a_819_n4851# a_287_4981# a_761_n5981#
+ a_1551_3763# a_n29_n5981# a_503_n6069# a_503_1239# a_n661_1327# a_n1393_n4851# a_n445_n6069#
+ a_287_1327# a_761_n2327# a_n661_n3545# a_n819_3763# a_187_3675# a_n29_n2327# a_1451_2457#
+ a_503_21# a_n919_n6069# a_1393_n5981# a_1135_n6069# a_n1551_n6069# a_n761_n4851#
+ a_n1451_4981# a_1393_n2327# a_187_n4851# a_n345_3763# a_n1451_1327# a_1451_n4851#
+ a_n187_109# a_n1609_3763# a_1235_2545# a_n603_4893# a_345_n6069# a_n287_n6069# a_1135_4893#
+ a_287_109# a_n1393_4893# a_819_n6069# a_n603_1239# a_129_n4763# a_1135_1239# a_761_2545#
+ a_n977_n3545# a_661_n4851# a_n287_3675# a_n1393_1239# a_n1393_n6069# a_661_4893#
+ a_919_4981# a_129_n1109# a_n1135_3763# a_n1135_n5981# a_661_1239# a_919_1327# a_n129_n3633#
+ a_1293_n4851# a_819_3675# a_n977_3763# a_n1609_n5981# a_n761_n6069# a_n1135_n2327#
+ a_1135_21# a_187_n6069# a_n503_n5981# a_603_n4763# a_n919_21# a_n1609_n2327# a_445_4981#
+ a_n1077_3675# a_n1235_n3633# a_1451_n6069# a_603_n1109# a_n503_n2327# a_n761_21#
+ a_n1753_n6203# a_n29_2545# a_445_1327# a_345_3675# a_n129_21# a_1235_n4763# a_977_n4851#
+ a_n603_n3633# a_n761_4893# a_1393_2545# a_n819_109# a_1293_4893# a_1235_n1109# a_661_n6069#
+ a_919_109# a_n761_1239# a_1293_1239# a_n919_3675# a_n345_n5981# a_n503_3763# a_445_n4763#
+ a_129_3763# a_n1077_n3633# a_1293_n6069# a_n1293_3763# a_n819_n5981# a_919_n4763#
+ a_445_n1109# a_n345_n2327# a_1077_4981# a_n1551_4893# a_n1451_n5981# a_1077_n4763#
+ a_977_3675# a_n187_2545# a_919_n1109# a_n819_n2327# a_503_n3633# a_n445_n3633# a_n661_109#
+ a_n445_3675# a_n1551_1239# a_1077_1327# a_n1393_21# a_29_n2415# a_n1451_n2327# a_1077_n1109#
+ a_761_109# a_n919_n3633# a_1135_n3633# a_n1551_n3633# a_977_n6069# a_819_21# a_n187_n5981#
+ a_287_n4763# a_661_21# a_29_2457# a_n187_n2327# a_1551_n4763# a_287_n1109# a_603_4981#
+ a_n1235_3675# a_n1293_n5981# a_345_n3633# a_1551_n1109# a_n287_n3633# a_603_1327#
+ a_n129_2457# a_n1293_n2327# a_503_3675# a_n661_3763# a_819_n3633# a_287_3763# a_n661_n5981#
+ a_761_n4763# a_1551_2545# a_n29_n4763# a_1451_4893# a_n1393_n3633# a_n661_n2327#
+ a_761_n1109# a_n819_2545# a_187_2457# a_1451_1239# a_n29_n1109# a_1393_n4763# a_n761_n3633#
+ a_29_n1197# a_n1451_3763# a_187_n3633# a_1393_n1109# a_1235_4981# a_1451_n3633#
+ a_n345_2545# a_n603_3675# a_n1609_2545# a_1235_1327# a_1293_21# a_1135_3675# a_761_4981#
+ a_n977_n5981# a_n1393_3675# a_129_n3545# a_761_1327# a_n977_n2327# a_661_n3633#
+ a_n287_2457# a_661_3675# a_919_3763# a_n287_21# a_n1135_2545# a_n1135_n4763# a_1293_n3633#
X0 a_n661_109# a_n761_21# a_n819_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X1 a_n187_n4763# a_n287_n4851# a_n345_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X2 a_1551_n5981# a_1451_n6069# a_1393_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X3 a_n29_n5981# a_n129_n6069# a_n187_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X4 a_129_n2327# a_29_n2415# a_n29_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X5 a_761_4981# a_661_4893# a_603_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X6 a_1393_2545# a_1293_2457# a_1235_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X7 a_n187_4981# a_n287_4893# a_n345_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X8 a_n1293_2545# a_n1393_2457# a_n1451_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X9 a_129_109# a_29_21# a_n29_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X10 a_445_n1109# a_345_n1197# a_287_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X11 a_287_3763# a_187_3675# a_129_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X12 a_n187_109# a_n287_21# a_n345_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X13 a_n187_n5981# a_n287_n6069# a_n345_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X14 a_129_n3545# a_29_n3633# a_n29_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X15 a_n1293_3763# a_n1393_3675# a_n1451_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X16 a_1393_3763# a_1293_3675# a_1235_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X17 a_n345_1327# a_n445_1239# a_n503_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X18 a_445_n2327# a_345_n2415# a_287_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X19 a_287_4981# a_187_4893# a_129_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X20 a_919_n1109# a_819_n1197# a_761_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X21 a_n819_109# a_n919_21# a_n977_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X22 a_129_n4763# a_29_n4851# a_n29_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X23 a_n1293_4981# a_n1393_4893# a_n1451_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X24 a_1393_4981# a_1293_4893# a_1235_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X25 a_129_1327# a_29_1239# a_n29_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X26 a_n345_109# a_n445_21# a_n503_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X27 a_n345_2545# a_n445_2457# a_n503_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X28 a_445_n3545# a_345_n3633# a_287_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X29 a_445_1327# a_345_1239# a_287_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X30 a_n1451_n1109# a_n1551_n1197# a_n1609_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X31 a_919_n2327# a_819_n2415# a_761_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X32 a_1077_n1109# a_977_n1197# a_919_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X33 a_129_n5981# a_29_n6069# a_n29_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X34 a_129_2545# a_29_2457# a_n29_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X35 a_n345_3763# a_n445_3675# a_n503_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X36 a_n1451_1327# a_n1551_1239# a_n1609_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X37 a_1551_1327# a_1451_1239# a_1393_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X38 a_445_n4763# a_345_n4851# a_287_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X39 a_n503_109# a_n603_21# a_n661_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X40 a_445_2545# a_345_2457# a_287_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X41 a_919_n3545# a_819_n3633# a_761_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X42 a_1077_n2327# a_977_n2415# a_919_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X43 a_n1451_n2327# a_n1551_n2415# a_n1609_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X44 a_n345_n1109# a_n445_n1197# a_n503_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X45 a_129_3763# a_29_3675# a_n29_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X46 a_1551_2545# a_1451_2457# a_1393_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X47 a_n345_4981# a_n445_4893# a_n503_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X48 a_n1451_2545# a_n1551_2457# a_n1609_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X49 a_445_n5981# a_345_n6069# a_287_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X50 a_n29_109# a_n129_21# a_n187_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X51 a_445_3763# a_345_3675# a_287_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X52 a_n977_1327# a_n1077_1239# a_n1135_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X53 a_919_n4763# a_819_n4851# a_761_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X54 a_1077_n3545# a_977_n3633# a_919_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X55 a_n1451_n3545# a_n1551_n3633# a_n1609_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X56 a_n345_n2327# a_n445_n2415# a_n503_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X57 a_129_4981# a_29_4893# a_n29_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X58 a_1551_3763# a_1451_3675# a_1393_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X59 a_1077_1327# a_977_1239# a_919_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X60 a_n1451_3763# a_n1551_3675# a_n1609_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X61 a_1393_109# a_1293_21# a_1235_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X62 a_n503_1327# a_n603_1239# a_n661_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X63 a_n819_n1109# a_n919_n1197# a_n977_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X64 a_445_4981# a_345_4893# a_287_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X65 a_n977_2545# a_n1077_2457# a_n1135_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X66 a_919_n5981# a_819_n6069# a_761_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X67 a_1077_n4763# a_977_n4851# a_919_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X68 a_n1451_n4763# a_n1551_n4851# a_n1609_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X69 a_1077_109# a_977_21# a_919_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X70 a_n977_n1109# a_n1077_n1197# a_n1135_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X71 a_n345_n3545# a_n445_n3633# a_n503_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X72 a_1551_4981# a_1451_4893# a_1393_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X73 a_1077_2545# a_977_2457# a_919_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X74 a_n1451_4981# a_n1551_4893# a_n1609_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X75 a_1235_n1109# a_1135_n1197# a_1077_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X76 a_n503_2545# a_n603_2457# a_n661_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X77 a_1551_109# a_1451_21# a_1393_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X78 a_n819_n2327# a_n919_n2415# a_n977_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X79 a_n977_3763# a_n1077_3675# a_n1135_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X80 a_1077_n5981# a_977_n6069# a_919_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X81 a_n1451_n5981# a_n1551_n6069# a_n1609_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X82 a_n29_1327# a_n129_1239# a_n187_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X83 a_603_1327# a_503_1239# a_445_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X84 a_n977_n2327# a_n1077_n2415# a_n1135_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X85 a_n345_n4763# a_n445_n4851# a_n503_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X86 a_1077_3763# a_977_3675# a_919_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X87 a_1235_n2327# a_1135_n2415# a_1077_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X88 a_1393_n1109# a_1293_n1197# a_1235_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X89 a_n503_3763# a_n603_3675# a_n661_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X90 a_761_109# a_661_21# a_603_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X91 a_n819_n3545# a_n919_n3633# a_n977_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X92 a_603_n1109# a_503_n1197# a_445_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X93 a_n977_4981# a_n1077_4893# a_n1135_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X94 a_n29_2545# a_n129_2457# a_n187_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X95 a_603_2545# a_503_2457# a_445_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X96 a_n977_n3545# a_n1077_n3633# a_n1135_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X97 a_n345_n5981# a_n445_n6069# a_n503_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X98 a_1077_4981# a_977_4893# a_919_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X99 a_1235_n3545# a_1135_n3633# a_1077_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X100 a_1393_n2327# a_1293_n2415# a_1235_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X101 a_n503_4981# a_n603_4893# a_n661_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X102 a_287_109# a_187_21# a_129_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X103 a_n819_n4763# a_n919_n4851# a_n977_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X104 a_603_n2327# a_503_n2415# a_445_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X105 a_761_n1109# a_661_n1197# a_603_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X106 a_1235_1327# a_1135_1239# a_1077_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X107 a_1235_109# a_1135_21# a_1077_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X108 a_n29_3763# a_n129_3675# a_n187_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X109 a_603_3763# a_503_3675# a_445_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X110 a_n1135_1327# a_n1235_1239# a_n1293_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X111 a_n977_n4763# a_n1077_n4851# a_n1135_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X112 a_1235_n4763# a_1135_n4851# a_1077_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X113 a_1393_n3545# a_1293_n3633# a_1235_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X114 a_919_109# a_819_21# a_761_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X115 a_n819_n5981# a_n919_n6069# a_n977_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X116 a_603_n3545# a_503_n3633# a_445_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X117 a_761_n2327# a_661_n2415# a_603_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X118 a_1235_2545# a_1135_2457# a_1077_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X119 a_445_109# a_345_21# a_287_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X120 a_n29_4981# a_n129_4893# a_n187_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X121 a_603_4981# a_503_4893# a_445_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X122 a_n1135_2545# a_n1235_2457# a_n1293_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X123 a_n977_n5981# a_n1077_n6069# a_n1135_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X124 a_1235_n5981# a_1135_n6069# a_1077_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X125 a_1393_n4763# a_1293_n4851# a_1235_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X126 a_761_n3545# a_661_n3633# a_603_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X127 a_603_n4763# a_503_n4851# a_445_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X128 a_1235_3763# a_1135_3675# a_1077_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X129 a_n1135_3763# a_n1235_3675# a_n1293_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X130 a_603_109# a_503_21# a_445_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X131 a_1393_n5981# a_1293_n6069# a_1235_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X132 a_n503_n1109# a_n603_n1197# a_n661_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X133 a_761_n4763# a_661_n4851# a_603_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X134 a_603_n5981# a_503_n6069# a_445_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X135 a_287_n1109# a_187_n1197# a_129_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X136 a_1235_4981# a_1135_4893# a_1077_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X137 a_n1135_4981# a_n1235_4893# a_n1293_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X138 a_n661_n1109# a_n761_n1197# a_n819_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X139 a_n503_n2327# a_n603_n2415# a_n661_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X140 a_761_n5981# a_661_n6069# a_603_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X141 a_287_n2327# a_187_n2415# a_129_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X142 a_n1135_n1109# a_n1235_n1197# a_n1293_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X143 a_n661_n2327# a_n761_n2415# a_n819_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X144 a_n1293_109# a_n1393_21# a_n1451_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X145 a_n503_n3545# a_n603_n3633# a_n661_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X146 a_n819_1327# a_n919_1239# a_n977_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X147 a_287_n3545# a_187_n3633# a_129_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X148 a_n1293_n1109# a_n1393_n1197# a_n1451_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X149 a_n661_1327# a_n761_1239# a_n819_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X150 a_n661_n3545# a_n761_n3633# a_n819_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X151 a_n1135_n2327# a_n1235_n2415# a_n1293_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X152 a_n503_n4763# a_n603_n4851# a_n661_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X153 a_n1451_109# a_n1551_21# a_n1609_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X154 a_1551_n1109# a_1451_n1197# a_1393_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X155 a_n29_n1109# a_n129_n1197# a_n187_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X156 a_n819_2545# a_n919_2457# a_n977_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X157 a_287_n4763# a_187_n4851# a_129_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X158 a_919_1327# a_819_1239# a_761_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X159 a_n1293_n2327# a_n1393_n2415# a_n1451_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X160 a_n661_2545# a_n761_2457# a_n819_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X161 a_n661_n4763# a_n761_n4851# a_n819_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X162 a_n1135_n3545# a_n1235_n3633# a_n1293_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X163 a_n503_n5981# a_n603_n6069# a_n661_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X164 a_n187_n1109# a_n287_n1197# a_n345_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X165 a_n819_3763# a_n919_3675# a_n977_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X166 a_n977_109# a_n1077_21# a_n1135_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X167 a_1551_n2327# a_1451_n2415# a_1393_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X168 a_n29_n2327# a_n129_n2415# a_n187_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X169 a_n187_1327# a_n287_1239# a_n345_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X170 a_761_1327# a_661_1239# a_603_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X171 a_287_n5981# a_187_n6069# a_129_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X172 a_919_2545# a_819_2457# a_761_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X173 a_n1293_n3545# a_n1393_n3633# a_n1451_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X174 a_n661_3763# a_n761_3675# a_n819_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X175 a_n661_n5981# a_n761_n6069# a_n819_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X176 a_n1135_n4763# a_n1235_n4851# a_n1293_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X177 a_n187_n2327# a_n287_n2415# a_n345_n2327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X178 a_n819_4981# a_n919_4893# a_n977_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X179 a_1551_n3545# a_1451_n3633# a_1393_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X180 a_n29_n3545# a_n129_n3633# a_n187_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X181 a_n187_2545# a_n287_2457# a_n345_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X182 a_761_2545# a_661_2457# a_603_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X183 a_n1135_109# a_n1235_21# a_n1293_109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X184 a_919_3763# a_819_3675# a_761_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X185 a_n1293_n4763# a_n1393_n4851# a_n1451_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X186 a_n661_4981# a_n761_4893# a_n819_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X187 a_287_1327# a_187_1239# a_129_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X188 a_n1135_n5981# a_n1235_n6069# a_n1293_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X189 a_n187_n3545# a_n287_n3633# a_n345_n3545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X190 a_1551_n4763# a_1451_n4851# a_1393_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X191 a_n29_n4763# a_n129_n4851# a_n187_n4763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X192 a_129_n1109# a_29_n1197# a_n29_n1109# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X193 a_761_3763# a_661_3675# a_603_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X194 a_1393_1327# a_1293_1239# a_1235_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X195 a_n187_3763# a_n287_3675# a_n345_3763# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X196 a_n1293_1327# a_n1393_1239# a_n1451_1327# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X197 a_919_4981# a_819_4893# a_761_4981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X198 a_n1293_n5981# a_n1393_n6069# a_n1451_n5981# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X199 a_287_2545# a_187_2457# a_129_2545# a_n1753_n6203# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_7EJ6Y6 a_n108_n250# w_n308_n547# a_50_n250# a_n50_n347#
X0 a_50_n250# a_n50_n347# a_n108_n250# w_n308_n547# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WSEQJ0 a_50_n200# a_n108_n200# a_n50_n288# a_n252_n422#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n252_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_L9TFKV a_n958_n300# a_n900_n388# a_n1092_n522#
+ a_900_n300#
X0 a_900_n300# a_n900_n388# a_n958_n300# a_n1092_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=9
.ends

.subckt sky130_am_ip__ldo_01v8 AVDD VOUT AVSS ENA VREF_EXT SEL_EXT DVDD DVSS
XXM56 vbias_p vy AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM67 vbias_n vbias_n vbias_n vbias_n AVSS AVSS vbias_n AVSS vbias_n vbias_n vbias_n
+ vbias_n AVSS AVSS AVSS vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM78 AVSS AVSS nena ena_3v3 sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0
XXM89 AVSS verr AVSS nena sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0
XXM46 vbias_p vx AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM57 vbias_c verr AVDD vy sky130_fd_pr__pfet_g5v0d10v5_KLAZY6__0
XXM68 AVDD vbias_c vbias_c AVDD sky130_fd_pr__pfet_g5v0d10v5_PC2PN5
XXM79 vbias_p vref_int AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
Xx1 ENA DVDD DVSS AVDD AVDD ena_3v3 AVDD DVSS DVSS sky130_fd_sc_hvl__lsbuflv2hv_1
XXM58 vbias_c m2_8539_n7649# AVDD vx sky130_fd_pr__pfet_g5v0d10v5_KLAZY6__0
XXM69 vbias_n vbias_n vbias_c vbias_n AVSS AVSS vbias_c AVSS vbias_c vbias_c vbias_c
+ vbias_n AVSS AVSS AVSS vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
Xx2 SEL_EXT DVDD DVSS AVDD AVDD sel_ext_3v3 AVDD DVSS DVSS sky130_fd_sc_hvl__lsbuflv2hv_1
XXM48 verr AVSS m2_8539_n7649# AVSS sky130_fd_pr__nfet_g5v0d10v5_69K6TN
XXM59 verr AVSS AVDD vpass sky130_fd_pr__pfet_g5v0d10v5_KLAZY6__0
XXR4 m1_5119_3142# m1_5119_2478# m1_5119_1150# m1_7519_2644# m1_7519_984# m1_7519_1980#
+ m1_5119_2146# m1_5119_3474# m1_7519_1648# m1_5119_1482# m1_7519_2976# m1_5119_2810#
+ vm m1_7519_2976# m1_5119_818# m1_5119_1814# m1_5119_1482# m1_7519_1316# m1_5119_3474#
+ m1_7519_3308# m1_5119_3142# m1_5119_2146# m1_7519_1648# m1_7519_2312# m1_7519_2644#
+ VOUT m1_5119_1150# AVSS m1_5119_2478# m1_7519_1316# m1_5119_2810# m1_7519_3308#
+ m1_7519_2312# m1_5119_818# m1_7519_1980# m1_5119_1814# m1_7519_984# sky130_fd_pr__res_xhigh_po_0p35_QZEXQH
XXR5 m1_5117_n1479# m1_5117_n2475# m1_7517_n4965# m1_5117_n4799# m1_7517_n981# m1_5117_n3803#
+ m1_5117_181# m1_7517_n1977# m1_7517_n3637# m1_7517_n2641# m1_7517_n4633# m1_5117_n815#
+ m1_7517_15# m1_5117_n2475# m1_5117_n5463# m1_5117_n151# m1_5117_n4467# m1_7517_n649#
+ m1_5117_n3471# m1_7517_n2973# m1_5117_n1147# vm m1_7517_n1645# m1_5117_181# m1_5117_n2143#
+ m1_7517_n3969# m1_7517_n4965# m1_5117_n815# m1_5117_n5131# m1_5117_n4135# m1_7517_n1977#
+ m1_5117_n2807# m1_7517_n981# m1_5117_n483# m1_7517_15# m1_7517_n3305# m1_5117_n3139#
+ m1_7517_n4301# m1_7517_n5297# m1_5117_n1479# m1_7517_n1645# m1_7517_n649# m1_7517_n4301#
+ m1_5117_n1811# m1_5117_n2807# m1_7517_n3305# m1_5117_n5463# m1_7517_n5297# m1_5117_n4467#
+ m1_7517_n2641# m1_5117_n151# m1_7517_n2309# m1_7517_n1313# m1_5117_n3471# m1_7517_n317#
+ m1_7517_n4633# m1_5117_n2143# m1_5117_n4799# m1_7517_n3637# AVSS AVSS m1_5117_n1147#
+ m1_5117_n1811# m1_5117_n5131# m1_7517_n1313# m1_5117_n3803# m1_7517_n2309# m1_5117_n483#
+ m1_5117_n4135# m1_7517_n3969# m1_7517_n317# m1_5117_n3139# m1_7517_n2973# sky130_fd_pr__res_xhigh_po_0p35_Z7JM9H
XXR6 AVSS m1_22164_n7435# AVSS m1_22164_n7435# m2_26640_n7437# sky130_fd_pr__res_xhigh_po_0p35_743D3R
XXC1[0] verr AVSS sky130_fd_pr__cap_mim_m3_1_MRZGNS
XXC1[1] verr AVSS sky130_fd_pr__cap_mim_m3_1_MRZGNS
XXC1[2] verr AVSS sky130_fd_pr__cap_mim_m3_1_MRZGNS
XXC3 AVSS vref sky130_fd_pr__cap_mim_m3_1_VCAG9S__0
XXM90 nena vdd_start AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_KLAZY6__0
XXM80 vref_int AVSS m1_12626_n9400# m1_10488_n8825# sky130_fd_pr__nfet_g5v0d10v5_PXBJUB
XXM70 AVSS vdd_start vbias_n vstart sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0
XXM81 vref_int AVSS vref_int m1_10488_n8825# sky130_fd_pr__nfet_g5v0d10v5_PXBJUB
XXM60 vbias_p vpass AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM71 m1_20910_n7332# vstart vstart AVDD sky130_fd_pr__pfet_g5v0d10v5_47NWVV
XXM82 vref_int AVSS m1_12626_n9400# AVSS sky130_fd_pr__nfet_g5v0d10v5_PXBJUB
XXM72 m1_20184_n7334# m1_20910_n7332# m1_20910_n7332# AVDD sky130_fd_pr__pfet_g5v0d10v5_47NWVV
XXM83 AVSS AVSS nsel_ext sel_ext_3v3 sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0
XXM61[0] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM61[1] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM61[2] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM61[3] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM61[4] vpass vpass AVDD AVDD VOUT vpass VOUT AVDD AVDD AVDD AVDD VOUT VOUT vpass
+ vpass VOUT VOUT AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass vpass AVDD VOUT
+ VOUT VOUT vpass VOUT AVDD VOUT AVDD AVDD vpass vpass VOUT VOUT vpass VOUT vpass
+ VOUT VOUT vpass vpass vpass vpass VOUT AVDD VOUT vpass vpass vpass vpass vpass VOUT
+ AVDD vpass vpass AVDD VOUT AVDD vpass AVDD vpass vpass vpass AVDD vpass VOUT AVDD
+ vpass vpass AVDD vpass vpass vpass AVDD AVDD VOUT AVDD VOUT AVDD vpass vpass vpass
+ vpass AVDD VOUT vpass VOUT vpass vpass vpass AVDD VOUT vpass vpass AVDD AVDD AVDD
+ vpass AVDD vpass vpass vpass AVDD VOUT vpass vpass VOUT AVDD vpass vpass VOUT vpass
+ VOUT AVDD vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass vpass VOUT AVDD VOUT
+ VOUT vpass vpass vpass vpass AVDD vpass AVDD AVDD vpass vpass AVDD VOUT AVDD VOUT
+ vpass VOUT vpass AVDD vpass vpass VOUT vpass AVDD vpass AVDD vpass vpass vpass vpass
+ vpass VOUT VOUT VOUT vpass vpass AVDD vpass AVDD VOUT vpass VOUT AVDD vpass VOUT
+ VOUT VOUT AVDD VOUT VOUT vpass AVDD vpass AVDD vpass vpass vpass VOUT vpass vpass
+ VOUT VOUT vpass vpass vpass vpass vpass vpass vpass AVDD AVDD vpass AVDD AVDD VOUT
+ VOUT vpass AVDD vpass vpass vpass vpass vpass AVDD vpass vpass AVDD vpass AVDD vpass
+ AVDD VOUT AVDD AVDD vpass vpass AVDD vpass vpass AVDD VOUT AVDD VOUT vpass AVDD
+ vpass vpass vpass VOUT vpass vpass vpass VOUT VOUT vpass AVDD VOUT vpass VOUT AVDD
+ AVDD vpass vpass vpass vpass AVDD vpass vpass vpass VOUT vpass VOUT AVDD vpass vpass
+ vpass vpass vpass AVDD VOUT VOUT VOUT vpass AVDD vpass vpass vpass AVDD AVDD vpass
+ VOUT vpass vpass VOUT AVDD vpass AVDD VOUT vpass vpass vpass AVDD VOUT vpass AVSS
+ AVDD VOUT vpass vpass AVDD vpass vpass vpass VOUT VOUT vpass AVDD vpass AVDD vpass
+ vpass vpass AVDD VOUT VOUT VOUT vpass vpass AVDD VOUT AVDD VOUT AVDD VOUT vpass
+ VOUT VOUT vpass VOUT AVDD VOUT vpass vpass AVDD vpass vpass VOUT vpass vpass VOUT
+ VOUT VOUT vpass vpass vpass vpass vpass VOUT AVDD vpass vpass VOUT AVDD AVDD AVDD
+ vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD vpass AVDD AVDD VOUT AVDD
+ AVDD vpass vpass AVDD VOUT VOUT vpass vpass AVDD VOUT vpass vpass VOUT vpass VOUT
+ AVDD vpass AVDD vpass AVDD AVDD vpass vpass VOUT AVDD vpass VOUT VOUT AVDD vpass
+ vpass vpass AVDD vpass VOUT VOUT vpass sky130_fd_pr__nfet_g5v0d10v5_YHRXVR
XXM62 vbias_p AVDD AVDD m1_19028_n7338# sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM73 AVDD m1_20184_n7334# m1_20184_n7334# AVDD sky130_fd_pr__pfet_g5v0d10v5_47NWVV
XXM84 AVDD AVDD nsel_ext sel_ext_3v3 sky130_fd_pr__pfet_g5v0d10v5_7EJ6Y6
Xsky130_fd_pr__pfet_g5v0d10v5_KLAZY6_0 ena_3v3 vbias_c AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_KLAZY6__0
XXM52 vy m2_6784_n8214# vm AVSS sky130_fd_pr__nfet_g5v0d10v5_WSEQJ0
XXM63 vbias_c m1_19028_n7338# AVDD vbias_p sky130_fd_pr__pfet_g5v0d10v5_KLAZY6__0
XXM74 vbias_n vbias_n vstart vbias_n AVSS AVSS vstart AVSS vstart vstart vstart vbias_n
+ AVSS AVSS AVSS vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM85 AVSS vbias_n AVSS nena sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0
XXM53 vx m2_6784_n8214# vref AVSS sky130_fd_pr__nfet_g5v0d10v5_WSEQJ0
XXM64 vbias_p AVDD AVDD m1_16878_n7330# sky130_fd_pr__pfet_g5v0d10v5_BWAZV5
XXM75 AVSS vref vref_int nsel_ext sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0
XXM54 AVSS vbias_n AVSS m2_6784_n8214# sky130_fd_pr__nfet_g5v0d10v5_L9TFKV
XXM65 vbias_c m1_16878_n7330# AVDD vbias_n sky130_fd_pr__pfet_g5v0d10v5_KLAZY6__0
XXM76 AVDD AVDD nena ena_3v3 sky130_fd_pr__pfet_g5v0d10v5_7EJ6Y6
XXM87 AVSS vpass AVSS nena sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0
XXM55 m2_8539_n7649# AVSS m2_8539_n7649# AVSS sky130_fd_pr__nfet_g5v0d10v5_69K6TN
XXM66[0] vbias_n vbias_n vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# vbias_p AVSS
+ vbias_p vbias_p vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# m2_26640_n7437#
+ vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM66[1] vbias_n vbias_n vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# vbias_p AVSS
+ vbias_p vbias_p vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# m2_26640_n7437#
+ vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM66[2] vbias_n vbias_n vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# vbias_p AVSS
+ vbias_p vbias_p vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# m2_26640_n7437#
+ vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM66[3] vbias_n vbias_n vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# vbias_p AVSS
+ vbias_p vbias_p vbias_p vbias_n m2_26640_n7437# m2_26640_n7437# m2_26640_n7437#
+ vbias_n sky130_fd_pr__nfet_g5v0d10v5_A2FZRM
XXM77 AVSS VREF_EXT vref sel_ext_3v3 sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N__0
XXM88 ena_3v3 vbias_p AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_KLAZY6__0
.ends

.subckt simple_switch_array_3 simplest_analog_switch_ena1v8_1[2]/in simplest_analog_switch_ena1v8_1[0]/on
+ simplest_analog_switch_ena1v8_1[0]/in simplest_analog_switch_ena1v8_1[1]/on simplest_analog_switch_ena1v8_1[1]/out
+ simplest_analog_switch_ena1v8_1[2]/on simplest_analog_switch_ena1v8_1[1]/in simplest_analog_switch_ena1v8_1[2]/avss
+ simplest_analog_switch_ena1v8_1[0]/out simplest_analog_switch_ena1v8_1[2]/out simplest_analog_switch_ena1v8_1[2]/dvdd
+ simplest_analog_switch_ena1v8_1[2]/avdd VSUBS
Xsimplest_analog_switch_ena1v8_1[0] simplest_analog_switch_ena1v8_1[2]/avdd simplest_analog_switch_ena1v8_1[2]/dvdd
+ simplest_analog_switch_ena1v8_1[2]/avss simplest_analog_switch_ena1v8_1[0]/on simplest_analog_switch_ena1v8_1[0]/out
+ VSUBS simplest_analog_switch_ena1v8_1[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1] simplest_analog_switch_ena1v8_1[2]/avdd simplest_analog_switch_ena1v8_1[2]/dvdd
+ simplest_analog_switch_ena1v8_1[2]/avss simplest_analog_switch_ena1v8_1[1]/on simplest_analog_switch_ena1v8_1[1]/out
+ VSUBS simplest_analog_switch_ena1v8_1[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[2] simplest_analog_switch_ena1v8_1[2]/avdd simplest_analog_switch_ena1v8_1[2]/dvdd
+ simplest_analog_switch_ena1v8_1[2]/avss simplest_analog_switch_ena1v8_1[2]/on simplest_analog_switch_ena1v8_1[2]/out
+ VSUBS simplest_analog_switch_ena1v8_1[2]/in simplest_analog_switch_ena1v8
.ends

.subckt sky130_fd_pr__nfet_01v8_QTPFY2 a_n29_n1250# a_n945_n1250# a_n429_n1338# a_945_n1338#
+ a_n487_n1250# a_n887_n1338# a_1803_n1250# a_487_n1338# a_1345_n1250# a_n1963_n1424#
+ a_n1403_n1250# a_n1803_n1338# a_429_n1250# a_n1861_n1250# a_887_n1250# a_n1345_n1338#
+ a_1403_n1338# a_29_n1338#
X0 a_n487_n1250# a_n887_n1338# a_n945_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=1.8125 pd=12.79 as=1.8125 ps=12.79 w=12.5 l=2
X1 a_n945_n1250# a_n1345_n1338# a_n1403_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=1.8125 pd=12.79 as=1.8125 ps=12.79 w=12.5 l=2
X2 a_887_n1250# a_487_n1338# a_429_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=1.8125 pd=12.79 as=1.8125 ps=12.79 w=12.5 l=2
X3 a_1803_n1250# a_1403_n1338# a_1345_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=3.625 pd=25.58 as=1.8125 ps=12.79 w=12.5 l=2
X4 a_1345_n1250# a_945_n1338# a_887_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=1.8125 pd=12.79 as=1.8125 ps=12.79 w=12.5 l=2
X5 a_n1403_n1250# a_n1803_n1338# a_n1861_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=1.8125 pd=12.79 as=3.625 ps=25.58 w=12.5 l=2
X6 a_n29_n1250# a_n429_n1338# a_n487_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=1.8125 pd=12.79 as=1.8125 ps=12.79 w=12.5 l=2
X7 a_429_n1250# a_29_n1338# a_n29_n1250# a_n1963_n1424# sky130_fd_pr__nfet_01v8 ad=1.8125 pd=12.79 as=1.8125 ps=12.79 w=12.5 l=2
.ends

.subckt sky130_fd_pr__nfet_01v8_QGRVRG a_n360_n674# a_200_n500# a_n258_n500# a_n200_n588#
X0 a_200_n500# a_n200_n588# a_n258_n500# a_n360_n674# sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=2
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_VCAG9S m3_n686_n540# c1_n646_n500#
X0 c1_n646_n500# m3_n686_n540# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
.ends

.subckt sky130_fd_pr__nfet_01v8_ME6MQD a_1000_n1000# a_n1160_n1174# a_n1000_n1088#
+ a_n1058_n1000#
X0 a_1000_n1000# a_n1000_n1088# a_n1058_n1000# a_n1160_n1174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=10
.ends

.subckt sky130_fd_pr__pfet_01v8_6H4ZLK a_n1000_n597# a_1000_n500# a_n1058_n500# w_n1196_n719#
X0 a_1000_n500# a_n1000_n597# a_n1058_n500# w_n1196_n719# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=10
.ends

.subckt sky130_fd_pr__nfet_01v8_D2R37Y a_1000_n500# a_n1058_n500# a_n1000_n588# a_n1160_n674#
X0 a_1000_n500# a_n1000_n588# a_n1058_n500# a_n1160_n674# sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=10
.ends

.subckt sky130_fd_pr__nfet_01v8_5TKQ2R a_500_n1000# a_n660_n1174# a_n500_n1088# a_n558_n1000#
X0 a_500_n1000# a_n500_n1088# a_n558_n1000# a_n660_n1174# sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=5
.ends

.subckt sbvfcm vdd pbias nbias vx vss XM7/w_n1196_n719# XM8/w_n1196_n719# VSUBS
Xsky130_fd_pr__nfet_01v8_QTPFY2_0 m1_5880_1010# m1_5880_1010# m1_5868_n3400# m1_5868_n3400#
+ vx m1_5868_n3400# m1_5880_1010# m1_5868_n3400# vx VSUBS vx m1_5868_n3400# vx m1_5880_1010#
+ m1_5880_1010# m1_5868_n3400# m1_5868_n3400# m1_5868_n3400# sky130_fd_pr__nfet_01v8_QTPFY2
XXM4 VSUBS m1_9368_n812# vss m1_5868_n3400# sky130_fd_pr__nfet_01v8_QGRVRG
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0 m1_9568_n2160# vdd sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXM5 pbias VSUBS nbias m1_5880_1010# sky130_fd_pr__nfet_01v8_ME6MQD
XXM6 m1_9368_n812# VSUBS nbias m1_5868_n3400# sky130_fd_pr__nfet_01v8_ME6MQD
XXM7 pbias pbias vdd XM7/w_n1196_n719# sky130_fd_pr__pfet_01v8_6H4ZLK
XXM8 pbias vdd m1_5868_n3400# XM8/w_n1196_n719# sky130_fd_pr__pfet_01v8_6H4ZLK
XXC1 m1_9568_n2160# vdd sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXM10 pbias vss m1_9568_n2160# VSUBS sky130_fd_pr__nfet_01v8_D2R37Y
XXM11 vss VSUBS m1_5868_n3400# m1_9568_n2160# sky130_fd_pr__nfet_01v8_5TKQ2R
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_H5FMR6 a_n199_n891# a_n69_n761# a_n69_329#
X0 a_n69_329# a_n69_n761# a_n199_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_H5TM75 a_n420_n761# a_n550_n891# a_n420_329#
+ a_48_n761# a_n186_n761# a_282_329# a_48_329# a_n186_329# a_282_n761#
X0 a_n420_329# a_n420_n761# a_n550_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X1 a_48_329# a_48_n761# a_n550_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X2 a_282_329# a_282_n761# a_n550_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X3 a_n186_329# a_n186_n761# a_n550_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
.ends

.subckt sky130_fd_pr__nfet_01v8_J222PV a_n429_n588# a_29_n588# a_n589_n674# a_n487_n500#
+ a_n29_n500# a_429_n500#
X0 a_n29_n500# a_n429_n588# a_n487_n500# a_n589_n674# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X1 a_429_n500# a_29_n588# a_n29_n500# a_n589_n674# sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_D5BT6X a_n420_n761# a_n654_329# a_n888_329#
+ a_n420_329# a_48_n761# a_n654_n761# a_n1018_n891# a_n888_n761# a_n186_n761# a_750_n761#
+ a_282_329# a_48_329# a_n186_329# a_282_n761# a_750_329# a_516_n761# a_516_329#
X0 a_n654_329# a_n654_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X1 a_n420_329# a_n420_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X2 a_48_329# a_48_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X3 a_282_329# a_282_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X4 a_n888_329# a_n888_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X5 a_750_329# a_750_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X6 a_516_329# a_516_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X7 a_n186_329# a_n186_n761# a_n1018_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_2G52HS a_48_n761# a_n186_n761# a_n316_n891#
+ a_48_329# a_n186_329#
X0 a_48_329# a_48_n761# a_n316_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
X1 a_n186_329# a_n186_n761# a_n316_n891# sky130_fd_pr__res_xhigh_po_0p69 l=3.45
.ends

.subckt trim_res A trim0 trim2 trim3 trim1 B VSUBS
Xsky130_fd_pr__res_xhigh_po_0p69_H5FMR6_0 VSUBS m1_835_n1590# B sky130_fd_pr__res_xhigh_po_0p69_H5FMR6
Xsky130_fd_pr__res_xhigh_po_0p69_H5TM75_0 m1_834_n3490# VSUBS m1_4520_n760# m1_4760_n1840#
+ m1_4760_n1840# m1_4980_n760# m1_4980_n760# m1_4520_n760# m1_1200_n3120# sky130_fd_pr__res_xhigh_po_0p69_H5TM75
XXM1 trim0 trim0 VSUBS B m1_835_n1590# B sky130_fd_pr__nfet_01v8_J222PV
XXM2 trim1 trim1 VSUBS m1_835_n1590# m1_834_n3490# m1_835_n1590# sky130_fd_pr__nfet_01v8_J222PV
XXM3 trim2 trim2 VSUBS m1_834_n3490# m1_1200_n3120# m1_834_n3490# sky130_fd_pr__nfet_01v8_J222PV
XXM4 trim3 trim3 VSUBS m1_1200_n3120# A m1_1200_n3120# sky130_fd_pr__nfet_01v8_J222PV
Xsky130_fd_pr__res_xhigh_po_0p69_D5BT6X_0 m1_4020_n3720# m1_3780_n2640# A m1_3780_n2640#
+ m1_4500_n3720# m1_3560_n3720# VSUBS m1_3560_n3720# m1_4020_n3720# m1_4960_n3720#
+ m1_4720_n2640# m1_4260_n2640# m1_4260_n2640# m1_4500_n3720# m1_1200_n3120# m1_4960_n3720#
+ m1_4720_n2640# sky130_fd_pr__res_xhigh_po_0p69_D5BT6X
Xsky130_fd_pr__res_xhigh_po_0p69_2G52HS_0 m1_834_n3490# m1_835_n1590# VSUBS m1_3920_n760#
+ m1_3920_n760# sky130_fd_pr__res_xhigh_po_0p69_2G52HS
.ends

.subckt sky130_fd_pr__nfet_01v8_QGMQL3 a_n158_n250# a_n100_n338# a_n260_n424# a_100_n250#
X0 a_100_n250# a_n100_n338# a_n158_n250# a_n260_n424# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_MMMA4V a_100_n500# a_n158_n500# a_n100_n588# a_n260_n674#
X0 a_100_n500# a_n100_n588# a_n158_n500# a_n260_n674# sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_HS3BL4 a_100_n800# a_n158_n800# a_n100_n888# a_n260_n974#
X0 a_100_n800# a_n100_n888# a_n158_n800# a_n260_n974# sky130_fd_pr__nfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_W2FWA4 a_n429_n588# a_29_n588# a_n589_n674# a_n487_n500#
+ a_n29_n500# a_429_n500#
X0 a_n29_n500# a_n429_n588# a_n487_n500# a_n589_n674# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=2
X1 a_429_n500# a_29_n588# a_n29_n500# a_n589_n674# sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=2
.ends

.subckt sky130_fd_pr__pfet_01v8_ST5LSM a_n1087_n2000# w_n1225_n2219# a_n1029_n2097#
+ a_n29_n2000# a_1029_n2000# a_29_n2097#
X0 a_n29_n2000# a_n1029_n2097# a_n1087_n2000# w_n1225_n2219# sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.29 as=5.8 ps=40.58 w=20 l=5
X1 a_1029_n2000# a_29_n2097# a_n29_n2000# w_n1225_n2219# sky130_fd_pr__pfet_01v8 ad=5.8 pd=40.58 as=2.9 ps=20.29 w=20 l=5
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_CXW7PW a_n487_n1000# a_429_n1000# a_29_n1088#
+ a_n621_n1222# a_n429_n1088# a_n29_n1000#
X0 a_429_n1000# a_29_n1088# a_n29_n1000# a_n621_n1222# sky130_fd_pr__nfet_05v0_nvt ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=2
X1 a_n29_n1000# a_n429_n1088# a_n487_n1000# a_n621_n1222# sky130_fd_pr__nfet_05v0_nvt ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=2
.ends

.subckt output_amp vo vp vn ibias vss vdd VSUBS
XXM1 ibias ibias VSUBS vss sky130_fd_pr__nfet_01v8_QGMQL3
XXM2 vss vcm ibias VSUBS sky130_fd_pr__nfet_01v8_MMMA4V
XXM3 vo vss ibias VSUBS sky130_fd_pr__nfet_01v8_HS3BL4
XXM4 vn vn VSUBS vcm m1_5267_n942# vcm sky130_fd_pr__nfet_01v8_W2FWA4
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[0] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[1] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[2] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[3] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
Xsky130_fd_pr__cap_mim_m3_1_VCAG9S_0[4] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXM5 vp vp VSUBS vcm m1_7167_n942# vcm sky130_fd_pr__nfet_01v8_J222PV
XXM6 m1_5168_2580# vdd m1_5168_2580# vdd sky130_fd_pr__pfet_01v8_6H4ZLK
XXM7 m1_5168_2580# vo_pre vdd vdd sky130_fd_pr__pfet_01v8_6H4ZLK
XXM8 vdd vdd vo_pre vo vdd vo_pre sky130_fd_pr__pfet_01v8_ST5LSM
XXM9 m1_5267_n942# m1_5267_n942# vn VSUBS vn m1_5168_2580# sky130_fd_pr__nfet_05v0_nvt_CXW7PW
XXC2[0] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXC2[1] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXC2[2] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXC2[3] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXC2[4] vo_pre vo sky130_fd_pr__cap_mim_m3_1_VCAG9S
XXM10 m1_7167_n942# m1_7167_n942# vp VSUBS vp vo_pre sky130_fd_pr__nfet_05v0_nvt_CXW7PW
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_E9MCU4 a_n433_n2363# a_n69_n2233# a_n69_1801#
+ a_165_1801# a_165_n2233# a_n303_n2233# a_n303_1801#
X0 a_n69_1801# a_n69_n2233# a_n433_n2363# sky130_fd_pr__res_xhigh_po_0p69 l=18.17
X1 a_165_1801# a_165_n2233# a_n433_n2363# sky130_fd_pr__res_xhigh_po_0p69 l=18.17
X2 a_n303_1801# a_n303_n2233# a_n433_n2363# sky130_fd_pr__res_xhigh_po_0p69 l=18.17
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_39QBTQ a_n69_844# a_n69_n1276# a_n199_n1406#
X0 a_n69_844# a_n69_n1276# a_n199_n1406# sky130_fd_pr__res_xhigh_po_0p69 l=8.6
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_NB3ZKH a_n420_1847# a_n186_n2279# a_n550_n2409#
+ a_48_1847# a_n186_1847# a_282_n2279# a_48_n2279# a_n420_n2279# a_282_1847#
X0 a_n186_1847# a_n186_n2279# a_n550_n2409# sky130_fd_pr__res_xhigh_po_0p69 l=18.63
X1 a_n420_1847# a_n420_n2279# a_n550_n2409# sky130_fd_pr__res_xhigh_po_0p69 l=18.63
X2 a_48_1847# a_48_n2279# a_n550_n2409# sky130_fd_pr__res_xhigh_po_0p69 l=18.63
X3 a_282_1847# a_282_n2279# a_n550_n2409# sky130_fd_pr__res_xhigh_po_0p69 l=18.63
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_GAZAU4 a_984_n2306# a_n186_1874# a_750_1874#
+ a_n1590_1874# a_984_1874# a_n1590_n2306# a_1218_n2306# a_282_n2306# a_n1720_n2436#
+ a_282_1874# a_48_n2306# a_n420_n2306# a_n1122_1874# a_1218_1874# a_750_n2306# a_516_1874#
+ a_n1356_1874# a_n1356_n2306# a_n420_1874# a_n888_n2306# a_516_n2306# a_48_1874#
+ a_n654_1874# a_n1122_n2306# a_n186_n2306# a_n888_1874# a_1452_n2306# a_1452_1874#
+ a_n654_n2306#
X0 a_282_1874# a_282_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X1 a_n654_1874# a_n654_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X2 a_n186_1874# a_n186_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X3 a_516_1874# a_516_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X4 a_n420_1874# a_n420_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X5 a_1452_1874# a_1452_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X6 a_n1590_1874# a_n1590_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X7 a_48_1874# a_48_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X8 a_984_1874# a_984_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X9 a_n1356_1874# a_n1356_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X10 a_1218_1874# a_1218_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X11 a_750_1874# a_750_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X12 a_n1122_1874# a_n1122_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
X13 a_n888_1874# a_n888_n2306# a_n1720_n2436# sky130_fd_pr__res_xhigh_po_0p69 l=18.9
.ends

.subckt sky130_fd_pr__nfet_01v8_2333C8 a_n2000_n338# a_n2160_n424# a_2000_n250# a_n2058_n250#
X0 a_2000_n250# a_n2000_n338# a_n2058_n250# a_n2160_n424# sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=20
.ends

.subckt sky130_fd_pr__nfet_01v8_Q33MQV a_1000_n200# a_n1058_n200# a_n1000_n288# a_n1160_n374#
X0 a_1000_n200# a_n1000_n288# a_n1058_n200# a_n1160_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=10
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
X0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 perim=2.64e+06 area=4.347e+11
.ends

.subckt sky130_fd_pr__pfet_01v8_B3G3L7 a_n29_n2618# a_n2029_21# a_29_21# w_n2225_n2837#
+ a_2029_118# a_2029_n2618# a_n2029_n2715# a_29_n2715# a_n2087_118# a_n29_118# a_n2087_n2618#
X0 a_2029_118# a_29_21# a_n29_118# w_n2225_n2837# sky130_fd_pr__pfet_01v8 ad=3.625 pd=25.58 as=1.8125 ps=12.79 w=12.5 l=10
X1 a_n29_118# a_n2029_21# a_n2087_118# w_n2225_n2837# sky130_fd_pr__pfet_01v8 ad=1.8125 pd=12.79 as=3.625 ps=25.58 w=12.5 l=10
X2 a_n29_n2618# a_n2029_n2715# a_n2087_n2618# w_n2225_n2837# sky130_fd_pr__pfet_01v8 ad=1.8125 pd=12.79 as=3.625 ps=25.58 w=12.5 l=10
X3 a_2029_n2618# a_29_n2715# a_n29_n2618# w_n2225_n2837# sky130_fd_pr__pfet_01v8 ad=3.625 pd=25.58 as=1.8125 ps=12.79 w=12.5 l=10
.ends

.subckt sky130_fd_pr__pfet_01v8_XPMKX6 a_30_n1000# a_n33_n1097# a_n88_n1000# w_n226_n1219#
X0 a_30_n1000# a_n33_n1097# a_n88_n1000# w_n226_n1219# sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.3
.ends

.subckt sky130_ak_ip__cmos_vref vbg avdd18 ena vbgsc vbgtg trim3 trim2 trim1 trim0
+ vptat dvdd dvss avss
Xsky130_fd_sc_hd__buf_1_4 trim1 dvss dvss dvdd dvdd trim1buf sky130_fd_sc_hd__buf_1
Xx1 avdd_ena pbias vref vptat avss avdd_ena avdd_ena avss sbvfcm
Xx3 x3/A trim0buf trim2buf trim3buf trim1buf avss avss trim_res
Xx2 vbg vref x2/vn x2/ibias avss avdd_ena avss output_amp
XR1 avss m1_9471_n10626# m1_9471_n10158# vbgtg m1_9471_n10626# m1_9471_n10158# vbg
+ sky130_fd_pr__res_xhigh_po_0p69_E9MCU4
XR2 vbgtg vbgsc avss sky130_fd_pr__res_xhigh_po_0p69_39QBTQ
XR3 vbgsc m1_9472_n11356# avss m1_13592_n11600# m1_13592_n11600# m1_9472_n11824# m1_9472_n11824#
+ m1_9472_n11356# x2/vn sky130_fd_pr__res_xhigh_po_0p69_NB3ZKH
XR4 m1_13651_n12750# m1_9472_n13920# m1_9472_n12984# m1_9472_n15324# m1_9472_n12984#
+ x3/A m1_13651_n12750# m1_13651_n13686# avss m1_9472_n13452# m1_13651_n13686# m1_13651_n14154#
+ m1_9472_n14856# m1_9472_n12516# m1_13651_n13218# m1_9472_n13452# m1_9472_n15324#
+ m1_13651_n15090# m1_9472_n14388# m1_13651_n14622# m1_13651_n13218# m1_9472_n13920#
+ m1_9472_n14388# m1_13651_n15090# m1_13651_n14154# m1_9472_n14856# x2/vn m1_9472_n12516#
+ m1_13651_n14622# sky130_fd_pr__res_xhigh_po_0p69_GAZAU4
XXM1 vref avss vptat avss sky130_fd_pr__nfet_01v8_2333C8
XXM2 vptat vref vref avss sky130_fd_pr__nfet_01v8_Q33MQV
Xsky130_fd_sc_hd__inv_2_0 ena dvss dvss dvdd dvdd sky130_fd_sc_hd__inv_2_0/Y sky130_fd_sc_hd__inv_2
XXM3 pbias x2/ibias avdd_ena avdd_ena sky130_fd_pr__pfet_01v8_6H4ZLK
Xsky130_fd_sc_hd__diode_2_0 trim2 dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
XXM9 vref pbias pbias avdd_ena avdd_ena avdd_ena pbias pbias avdd_ena vref avdd_ena
+ sky130_fd_pr__pfet_01v8_B3G3L7
Xsky130_fd_sc_hd__diode_2_1 ena dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_2 trim3 dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_3 trim1 dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__decap_6_0 dvss dvss dvdd dvdd sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__diode_2_4 trim0 dvss dvss dvdd dvdd sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__buf_1_0 trim0 dvss dvss dvdd dvdd trim0buf sky130_fd_sc_hd__buf_1
XXM20 avdd_ena sky130_fd_sc_hd__inv_2_0/Y avdd18 dvdd sky130_fd_pr__pfet_01v8_XPMKX6
Xsky130_fd_sc_hd__buf_1_2 trim3 dvss dvss dvdd dvdd trim3buf sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_3 trim2 dvss dvss dvdd dvdd trim2buf sky130_fd_sc_hd__buf_1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N a_n252_n322# a_50_n100# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n252_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_VHBZVD a_n400_n197# a_400_n100# w_n658_n397#
+ a_n458_n100#
X0 a_400_n100# a_n400_n197# a_n458_n100# w_n658_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3 a_50_n400# a_n247_n622# a_n108_n400# a_n50_n488#
X0 a_50_n400# a_n50_n488# a_n108_n400# a_n247_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLNSY6 a_n29_n100# w_n387_n397# a_n187_n100#
+ a_29_n197# a_n129_n197# a_129_n100#
X0 a_129_n100# a_29_n197# a_n29_n100# w_n387_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n197# a_n187_n100# w_n387_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLAZY6 a_n50_n197# a_50_n100# w_n308_n397# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n308_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_T4TNG7 a_n100_n597# a_n100_21# a_100_109# a_100_n509#
+ a_n158_n509# a_n158_109# a_n297_n731#
X0 a_100_n509# a_n100_n597# a_n158_n509# a_n297_n731# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X1 a_100_109# a_n100_21# a_n158_109# a_n297_n731# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_SALWK2 a_n88_n400# a_n33_n488# a_n190_n574# a_30_n400#
X0 a_30_n400# a_n33_n488# a_n88_n400# a_n190_n574# sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.3
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGK6VM a_n100_n297# a_100_n200# w_n358_n497#
+ a_n158_n200#
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n358_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_FVGVKR a_n284_684# a_214_n1116# a_n118_684#
+ a_48_n1116# a_n284_n1116# a_n414_n1246# a_n118_n1116# a_48_684# a_214_684#
X0 a_214_684# a_214_n1116# a_n414_n1246# sky130_fd_pr__res_xhigh_po_0p35 l=7
X1 a_n284_684# a_n284_n1116# a_n414_n1246# sky130_fd_pr__res_xhigh_po_0p35 l=7
X2 a_48_684# a_48_n1116# a_n414_n1246# sky130_fd_pr__res_xhigh_po_0p35 l=7
X3 a_n118_684# a_n118_n1116# a_n414_n1246# sky130_fd_pr__res_xhigh_po_0p35 l=7
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KL3SY6 a_n50_n497# a_50_n400# w_n308_n697# a_n108_n400#
X0 a_50_n400# a_n50_n497# a_n108_n400# w_n308_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_B8TQK3 a_n100_n597# a_n100_21# a_n260_n683# a_100_109#
+ a_100_n509# a_n158_n509# a_n158_109#
X0 a_100_n509# a_n100_n597# a_n158_n509# a_n260_n683# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X1 a_100_109# a_n100_21# a_n158_109# a_n260_n683# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt comparator_final Vinn Vinp RST AVDD DVDD ibn180n vo VSS
XXM12 VSS m1_9711_n5360# VSS vo1 sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM23 m2_26_n3922# m2_26_n3922# AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_VHBZVD
XXM14 vo1 VSS VSS vo sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3
XXM13 m1_9711_n5360# DVDD DVDD vo1 vo1 DVDD sky130_fd_pr__pfet_g5v0d10v5_KLNSY6
XXM24 m2_26_n3922# vbn AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_VHBZVD
XXM15 vo vo1 li_9669_n4446# li_9669_n4446# sky130_fd_pr__pfet_g5v0d10v5_KLAZY6
XXM26 vbn vbn VSS VSS vbn ibn180n VSS sky130_fd_pr__nfet_g5v0d10v5_T4TNG7
XXM16 VSS RST VSS m1_9711_n5360# sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N
XXM27 m2_26_n3922# VSS vbn m2_n888_n4722# sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3
XXM17 RST DVDD DVDD m1_9711_n5360# m1_9711_n5360# DVDD sky130_fd_pr__pfet_g5v0d10v5_KLNSY6
XXM28 VSS vbn VSS m2_n888_n4722# sky130_fd_pr__nfet_01v8_SALWK2
XXM19 li_9669_n4446# li_9669_n4446# AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_FGK6VM
XXR12 m1_2193_n3581# VSS m1_2193_n3581# m1_2360_n5380# m2_1724_n5235# VSS m1_2360_n5380#
+ m1_2525_n3581# m1_2525_n3581# sky130_fd_pr__res_xhigh_po_0p35_FVGVKR
XXM1 vbn vbn VS VS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_T4TNG7
XXM2 m1_7183_n5366# vt AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_KL3SY6
XXM3 m1_7183_n5366# m1_7183_n5366# AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_KL3SY6
XXM4 m1_7183_n5366# VSS m2_6521_n3805# AVDD sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3
XXM5 m1_n1718_n3574# m1_n1718_n3574# AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_VHBZVD
XXM6 vbn vbn VSS VSS vo vo VSS sky130_fd_pr__nfet_g5v0d10v5_T4TNG7
XXM7 vt AVDD AVDD vo sky130_fd_pr__pfet_g5v0d10v5_KL3SY6
XXM8 vt VSS m1_5358_n4724# AVDD sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3
Xsky130_fd_pr__nfet_01v8_B8TQK3_0 Vinn VSS VSS VSS VS m1_5358_n4724# VSS sky130_fd_pr__nfet_01v8_B8TQK3
Xsky130_fd_pr__nfet_01v8_B8TQK3_1 Vinn Vinn VSS VS VS m1_5358_n4724# m1_5358_n4724#
+ sky130_fd_pr__nfet_01v8_B8TQK3
Xsky130_fd_pr__nfet_01v8_B8TQK3_2 Vinn Vinn VSS VS VS m1_5358_n4724# m1_5358_n4724#
+ sky130_fd_pr__nfet_01v8_B8TQK3
Xsky130_fd_pr__nfet_01v8_B8TQK3_3 Vinn Vinn VSS VS VS m1_5358_n4724# m1_5358_n4724#
+ sky130_fd_pr__nfet_01v8_B8TQK3
Xsky130_fd_pr__nfet_g5v0d10v5_T4TNG7_0 vbn vbn m2_1724_n5235# m2_1724_n5235# m2_26_n3922#
+ m2_26_n3922# VSS sky130_fd_pr__nfet_g5v0d10v5_T4TNG7
XXM20 m2_n888_n4722# m2_n888_n4722# AVDD m1_n1844_n4683# sky130_fd_pr__pfet_g5v0d10v5_VHBZVD
XXM10 Vinp Vinp VSS m2_6521_n3805# m2_6521_n3805# VS VS sky130_fd_pr__nfet_01v8_B8TQK3
XXM11 m1_n1844_n4683# m1_n1718_n3574# AVDD m1_n1844_n4683# sky130_fd_pr__pfet_g5v0d10v5_VHBZVD
.ends

.subckt sky130_fd_pr__pfet_01v8_GHZ9W9 a_n29_n100# a_89_n100# a_26_n197# w_n285_n319#
+ a_n92_n197# a_n147_n100#
X0 a_n29_n100# a_n92_n197# a_n147_n100# w_n285_n319# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X1 a_89_n100# a_26_n197# a_n29_n100# w_n285_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
.ends

.subckt sky130_fd_pr__pfet_01v8_XPC8Y6 a_n29_n100# a_n187_n100# a_29_n197# a_n129_n197#
+ a_129_n100# w_n325_n319#
X0 a_129_n100# a_29_n197# a_n29_n100# w_n325_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n197# a_n187_n100# w_n325_n319# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_L9ESAD a_n175_n224# a_n73_n50# a_n33_n154# a_15_n50#
X0 a_15_n50# a_n33_n154# a_n73_n50# a_n175_n224# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_2V27AY m4_200_n17880# c2_280_n17800# c2_n4018_n17800#
+ m4_n4098_n17880#
X0 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X1 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X2 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X3 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X4 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X5 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X6 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X7 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X8 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X9 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X10 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X11 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X12 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X13 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X14 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X15 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X16 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X17 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X18 c2_280_n17800# m4_200_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
X19 c2_n4018_n17800# m4_n4098_n17880# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
.ends

.subckt sky130_fd_pr__nfet_01v8_PR763Z a_591_n50# a_1071_n50# a_207_n50# a_n465_n50#
+ a_n207_n76# a_n945_n50# a_783_n50# a_1263_n50# a_n177_n50# a_n1299_72# a_n1427_n224#
+ a_n657_n50# a_n1137_n50# a_n1325_n50# a_495_n50# a_111_n50# a_975_n50# a_n369_n50#
+ a_n975_n76# a_n849_n50# a_1167_n50# a_687_n50# a_303_n50# a_n561_n50# a_n1041_n50#
+ a_n1167_n76# a_n81_n50# a_399_n50# a_879_n50# a_n273_n50# a_15_n50# a_n753_n50#
+ a_n1233_n50#
X0 a_15_n50# a_n207_n76# a_n81_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X1 a_111_n50# a_n207_n76# a_15_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X2 a_n273_n50# a_n975_n76# a_n369_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X3 a_n81_n50# a_n207_n76# a_n177_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X4 a_n177_n50# a_n207_n76# a_n273_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X5 a_303_n50# a_n207_n76# a_207_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X6 a_591_n50# a_n207_n76# a_495_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X7 a_207_n50# a_n207_n76# a_111_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X8 a_399_n50# a_n207_n76# a_303_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X9 a_495_n50# a_n207_n76# a_399_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X10 a_687_n50# a_n207_n76# a_591_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X11 a_783_n50# a_n207_n76# a_687_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X12 a_975_n50# a_n207_n76# a_879_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X13 a_n1041_n50# a_n1167_n76# a_n1137_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X14 a_879_n50# a_n207_n76# a_783_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X15 a_n1233_n50# a_n1299_72# a_n1325_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.155 ps=1.62 w=0.5 l=0.15
X16 a_n1137_n50# a_n1167_n76# a_n1233_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X17 a_n561_n50# a_n975_n76# a_n657_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X18 a_1071_n50# a_n207_n76# a_975_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X19 a_1167_n50# a_n207_n76# a_1071_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X20 a_1263_n50# a_n207_n76# a_1167_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.155 pd=1.62 as=0.0825 ps=0.83 w=0.5 l=0.15
X21 a_n945_n50# a_n975_n76# a_n1041_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X22 a_n849_n50# a_n975_n76# a_n945_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X23 a_n753_n50# a_n975_n76# a_n849_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X24 a_n657_n50# a_n975_n76# a_n753_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X25 a_n465_n50# a_n975_n76# a_n561_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
X26 a_n369_n50# a_n975_n76# a_n465_n50# a_n1427_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.0825 ps=0.83 w=0.5 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_DD63S8 a_n465_n202# a_n945_18# a_1167_n202# a_n81_18#
+ a_n273_18# a_15_n202# a_n561_n202# a_975_18# a_n177_n202# a_303_18# a_1263_n202#
+ a_879_n202# a_111_n202# a_n1041_18# a_n975_n299# a_n273_n202# a_n1137_n202# a_n849_18#
+ a_975_n202# a_n561_18# a_1071_18# a_879_18# a_n177_18# a_n1233_n202# a_207_18# a_591_18#
+ a_1071_n202# a_687_n202# a_15_18# a_n465_18# a_783_n202# a_399_n202# a_n81_n202#
+ a_n849_n202# w_n1463_n397# a_495_18# a_n1233_18# a_n1041_n202# a_n1299_n299# a_495_n202#
+ a_n945_n202# a_n753_18# a_1263_18# a_n369_18# a_783_18# a_n1137_18# a_n207_n299#
+ a_591_n202# a_n657_n202# a_399_18# a_111_18# a_207_n202# a_n1167_n299# a_n753_n202#
+ a_n1325_n202# a_1167_18# a_n657_18# a_n369_n202# a_n1325_18# a_303_n202# a_687_18#
X0 a_n1233_n202# a_n1299_n299# a_n1325_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X1 a_591_n202# a_n207_n299# a_495_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X2 a_n657_18# a_n975_n299# a_n753_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X3 a_975_18# a_n207_n299# a_879_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X4 a_1263_18# a_n207_n299# a_1167_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X5 a_n849_n202# a_n975_n299# a_n945_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X6 a_n945_18# a_n975_n299# a_n1041_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X7 a_879_18# a_n207_n299# a_783_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X8 a_n177_n202# a_n207_n299# a_n273_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X9 a_207_n202# a_n207_n299# a_111_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X10 a_1167_18# a_n207_n299# a_1071_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X11 a_n1137_n202# a_n1167_n299# a_n1233_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X12 a_495_n202# a_n207_n299# a_399_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X13 a_n849_18# a_n975_n299# a_n945_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X14 a_n81_18# a_n207_n299# a_n177_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X15 a_n561_n202# a_n975_n299# a_n657_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X16 a_111_n202# a_n207_n299# a_15_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X17 a_783_n202# a_n207_n299# a_687_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X18 a_1071_n202# a_n207_n299# a_975_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X19 a_303_18# a_n207_n299# a_207_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X20 a_399_n202# a_n207_n299# a_303_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X21 a_n1041_18# a_n1167_n299# a_n1137_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X22 a_n273_18# a_n975_n299# a_n369_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X23 a_111_18# a_n207_n299# a_15_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X24 a_n465_n202# a_n975_n299# a_n561_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X25 a_687_n202# a_n207_n299# a_591_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X26 a_207_18# a_n207_n299# a_111_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X27 a_591_18# a_n207_n299# a_495_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X28 a_n753_n202# a_n975_n299# a_n849_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X29 a_975_n202# a_n207_n299# a_879_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X30 a_n177_18# a_n207_n299# a_n273_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X31 a_15_18# a_n207_n299# a_n81_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X32 a_n81_n202# a_n207_n299# a_n177_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X33 a_1263_n202# a_n207_n299# a_1167_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X34 a_n561_18# a_n975_n299# a_n657_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X35 a_495_18# a_n207_n299# a_399_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X36 a_15_n202# a_n207_n299# a_n81_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X37 a_n1233_18# a_n1299_n299# a_n1325_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X38 a_n1041_n202# a_n1167_n299# a_n1137_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X39 a_n369_n202# a_n975_n299# a_n465_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X40 a_n465_18# a_n975_n299# a_n561_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X41 a_399_18# a_n207_n299# a_303_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X42 a_n657_n202# a_n975_n299# a_n753_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X43 a_n1137_18# a_n1167_n299# a_n1233_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X44 a_783_18# a_n207_n299# a_687_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X45 a_879_n202# a_n207_n299# a_783_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X46 a_1071_18# a_n207_n299# a_975_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X47 a_n945_n202# a_n975_n299# a_n1041_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X48 a_1167_n202# a_n207_n299# a_1071_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X49 a_n753_18# a_n975_n299# a_n849_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X50 a_n369_18# a_n975_n299# a_n465_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X51 a_303_n202# a_n207_n299# a_207_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X52 a_687_18# a_n207_n299# a_591_18# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
X53 a_n273_n202# a_n975_n299# a_n369_n202# w_n1463_n397# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.1155 ps=1.03 w=0.7 l=0.15
.ends

.subckt por_output_buffer w_33421_n285686# m2_34641_n286220# VSUBS m1_33354_n286009#
XXM53 m2_34641_n286220# VSUBS m2_34641_n286220# VSUBS m2_33873_n286220# m2_33873_n286220#
+ m2_34641_n286220# VSUBS m2_34641_n286220# m1_33354_n286009# VSUBS VSUBS m2_33681_n286220#
+ m2_33489_n286220# VSUBS VSUBS m2_34641_n286220# m2_33873_n286220# m2_33681_n286220#
+ VSUBS m2_34641_n286220# VSUBS VSUBS m2_33873_n286220# VSUBS m2_33489_n286220# VSUBS
+ m2_34641_n286220# VSUBS VSUBS m2_34641_n286220# m2_33873_n286220# VSUBS sky130_fd_pr__nfet_01v8_PR763Z
XXM54 w_33421_n285686# m2_33873_n286220# m2_34641_n286220# w_33421_n285686# w_33421_n285686#
+ m2_34641_n286220# m2_33873_n286220# m2_34641_n286220# m2_34641_n286220# w_33421_n285686#
+ w_33421_n285686# w_33421_n285686# w_33421_n285686# w_33421_n285686# m2_33681_n286220#
+ w_33421_n285686# m2_33681_n286220# w_33421_n285686# m2_34641_n286220# m2_33873_n286220#
+ w_33421_n285686# w_33421_n285686# m2_34641_n286220# w_33421_n285686# m2_34641_n286220#
+ m2_34641_n286220# w_33421_n285686# w_33421_n285686# m2_34641_n286220# w_33421_n285686#
+ m2_34641_n286220# m2_34641_n286220# w_33421_n285686# w_33421_n285686# w_33421_n285686#
+ w_33421_n285686# w_33421_n285686# w_33421_n285686# m1_33354_n286009# w_33421_n285686#
+ m2_33873_n286220# m2_33873_n286220# w_33421_n285686# m2_33873_n286220# m2_34641_n286220#
+ m2_33681_n286220# m2_33873_n286220# m2_34641_n286220# w_33421_n285686# m2_34641_n286220#
+ w_33421_n285686# m2_34641_n286220# m2_33489_n286220# m2_33873_n286220# m2_33489_n286220#
+ m2_34641_n286220# w_33421_n285686# m2_33873_n286220# m2_33489_n286220# w_33421_n285686#
+ w_33421_n285686# sky130_fd_pr__pfet_01v8_DD63S8
.ends

.subckt sky130_fd_pr__nfet_01v8_G7LLWL a_n29_n50# a_26_n154# a_n249_n224# a_n147_n50#
+ a_89_n50# a_n92_n154#
X0 a_89_n50# a_26_n154# a_n29_n50# a_n249_n224# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.3
X1 a_n29_n50# a_n92_n154# a_n147_n50# a_n249_n224# sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.3
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_PQJ659 a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__pfet_01v8_U6B66J a_n73_118# a_n33_21# w_n211_n477# a_n73_n258#
+ a_15_118# a_n33_n355# a_15_n258#
X0 a_15_118# a_n33_21# a_n73_118# w_n211_n477# sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.98 as=0.203 ps=1.98 w=0.7 l=0.15
X1 a_15_n258# a_n33_n355# a_n73_n258# w_n211_n477# sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.98 as=0.203 ps=1.98 w=0.7 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_SKYQWJ a_n88_n318# a_30_118# a_n33_n415# a_n33_21#
+ a_n88_118# a_30_n318# w_n226_n537#
X0 a_30_n318# a_n33_n415# a_n88_n318# w_n226_n537# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X1 a_30_118# a_n33_21# a_n88_118# w_n226_n537# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLZS5A a_n683_n200# a_n189_n297# a_29_n297# a_189_n200#
+ a_n901_n200# a_247_n297# a_n407_n297# a_465_n297# a_407_n200# a_n625_n297# a_683_n297#
+ a_625_n200# a_n843_n297# w_n1101_n497# a_843_n200# a_n29_n200# a_n247_n200# a_n465_n200#
X0 a_n247_n200# a_n407_n297# a_n465_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_843_n200# a_683_n297# a_625_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X2 a_407_n200# a_247_n297# a_189_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X3 a_189_n200# a_29_n297# a_n29_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n465_n200# a_n625_n297# a_n683_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_625_n200# a_465_n297# a_407_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_n29_n200# a_n189_n297# a_n247_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X7 a_n683_n200# a_n843_n297# a_n901_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__nfet_01v8_5QNSAB a_n33_n50# a_n227_n224# a_63_n50# a_n125_n50#
+ a_n81_n154#
X0 a_n33_n50# a_n81_n154# a_n125_n50# a_n227_n224# sky130_fd_pr__nfet_01v8 ad=0.0825 pd=0.83 as=0.155 ps=1.62 w=0.5 l=0.15
X1 a_63_n50# a_n81_n154# a_n33_n50# a_n227_n224# sky130_fd_pr__nfet_01v8 ad=0.155 pd=1.62 as=0.0825 ps=0.83 w=0.5 l=0.15
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WSE8X6 a_n331_n402# a_29_n268# a_n29_n180# a_n129_n268#
+ a_n187_n180# a_129_n180#
X0 a_129_n180# a_29_n268# a_n29_n180# a_n331_n402# sky130_fd_pr__nfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.261 ps=2.09 w=1.8 l=0.5
X1 a_n29_n180# a_n129_n268# a_n187_n180# a_n331_n402# sky130_fd_pr__nfet_g5v0d10v5 ad=0.261 pd=2.09 as=0.522 ps=4.18 w=1.8 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_PHU9Y6 a_129_n290# a_29_n387# a_n129_n387# a_n29_n290#
+ a_n187_n290# w_n387_n587#
X0 a_129_n290# a_29_n387# a_n29_n290# w_n387_n587# sky130_fd_pr__pfet_g5v0d10v5 ad=0.841 pd=6.38 as=0.4205 ps=3.19 w=2.9 l=0.5
X1 a_n29_n290# a_n129_n387# a_n187_n290# w_n387_n587# sky130_fd_pr__pfet_g5v0d10v5 ad=0.4205 pd=3.19 as=0.841 ps=6.38 w=2.9 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_X6X8XQ a_n81_n167# a_n33_n70# a_63_n70# a_n125_n70#
+ w_n263_n289#
X0 a_n33_n70# a_n81_n167# a_n125_n70# w_n263_n289# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X1 a_63_n70# a_n81_n167# a_n33_n70# w_n263_n289# sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_N5F8XL a_n108_n180# a_n242_n402# a_n50_n268#
+ a_50_n180#
X0 a_50_n180# a_n50_n268# a_n108_n180# a_n242_n402# sky130_fd_pr__nfet_g5v0d10v5 ad=0.522 pd=4.18 as=0.522 ps=4.18 w=1.8 l=0.5
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_FJFAMD m3_n386_n240# c1_n346_n200#
X0 c1_n346_n200# m3_n386_n240# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt levelShifter ain aout VCCL VSS VCCH
Xsky130_fd_pr__nfet_g5v0d10v5_WSE8X6_0 VSS S1B VSS S1B m2_2125_n529# m2_2125_n529#
+ sky130_fd_pr__nfet_g5v0d10v5_WSE8X6
XXM12 VSS S1 VSS S1 m1_2633_n381# m1_2633_n381# sky130_fd_pr__nfet_g5v0d10v5_WSE8X6
XXM13 m2_2125_n529# m1_2633_n381# m1_2633_n381# VCCH m2_2125_n529# VCCH sky130_fd_pr__pfet_g5v0d10v5_PHU9Y6
XXM1 ain VCCL S1 S1 VCCL sky130_fd_pr__pfet_01v8_X6X8XQ
XXM2 m1_2633_n381# m2_2125_n529# m2_2125_n529# VCCH m1_2633_n381# VCCH sky130_fd_pr__pfet_g5v0d10v5_PHU9Y6
XXM4 VSS VSS S1 S1B sky130_fd_pr__nfet_01v8_L9ESAD
XXM5 S1 VCCL S1B S1B VCCL sky130_fd_pr__pfet_01v8_X6X8XQ
XXM6 VSS VSS ain S1 sky130_fd_pr__nfet_01v8_L9ESAD
XXM7 aout VSS m2_2125_n529# VSS sky130_fd_pr__nfet_g5v0d10v5_N5F8XL
XXM8 aout m2_2125_n529# m2_2125_n529# VCCH aout VCCH sky130_fd_pr__pfet_g5v0d10v5_PHU9Y6
Xsky130_fd_pr__cap_mim_m3_1_FJFAMD_0 m2_2125_n529# VCCH sky130_fd_pr__cap_mim_m3_1_FJFAMD
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_69TNYL a_100_n100# a_n292_n322# a_n158_n100#
+ a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n292_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ESEQJ8 a_n282_n422# a_80_n200# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n282_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_TBT74C c1_n1746_n1600# m3_n1786_n1640#
X0 c1_n1746_n1600# m3_n1786_n1640# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_SYBQJL a_n792_n200# a_298_n200# a_516_n200# a_734_n200#
+ a_n926_n422# a_138_n288# a_n298_n288# a_80_n200# a_356_n288# a_n516_n288# a_574_n288#
+ a_n734_n288# a_n138_n200# a_n356_n200# a_n574_n200# a_n80_n288#
X0 a_n574_n200# a_n734_n288# a_n792_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X1 a_734_n200# a_574_n288# a_516_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X2 a_298_n200# a_138_n288# a_80_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X3 a_n138_n200# a_n298_n288# a_n356_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n356_n200# a_n516_n288# a_n574_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_516_n200# a_356_n288# a_298_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_80_n200# a_n80_n288# a_n138_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_KB5CJD m3_n1186_n1040# c1_n1146_n1000#
X0 c1_n1146_n1000# m3_n1186_n1040# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CAF9E7 a_29_n347# a_n129_n347# a_n29_n250# a_n187_n250#
+ w_n387_n547# a_129_n250#
X0 a_129_n250# a_29_n347# a_n29_n250# w_n387_n547# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=0.5
X1 a_n29_n250# a_n129_n347# a_n187_n250# w_n387_n547# sky130_fd_pr__pfet_g5v0d10v5 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_X6E435 a_n29_n100# a_n187_n100# a_129_n100# a_n331_n322#
+ a_29_n188# a_n129_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n331_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n188# a_n187_n100# a_n331_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_sc_hvl__inv_16 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X3 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X4 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X5 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X6 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X7 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X8 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X9 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X10 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X11 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X12 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X13 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X14 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X15 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X16 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X17 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X18 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X19 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X20 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X21 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.2025 pd=2.04 as=0.105 ps=1.03 w=0.75 l=0.5
X22 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X23 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X24 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X25 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X26 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X27 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X28 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X29 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X30 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X31 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt por_output_driver_h sky130_fd_sc_hvl__inv_16_0/VPWR sky130_fd_sc_hvl__inv_16_0/Y
+ sky130_fd_sc_hvl__inv_16_1/VPB sky130_fd_sc_hvl__inv_16_0/VGND sky130_fd_sc_hvl__inv_16_1/VPWR
+ m2_26866_n292108# m2_26862_n291518# sky130_fd_sc_hvl__inv_16_1/VGND sky130_fd_sc_hvl__inv_16_1/Y
+ VSUBS
Xsky130_fd_pr__pfet_g5v0d10v5_CAF9E7_0 m2_26960_n292468# m2_26960_n292468# m2_27646_n292468#
+ m2_26862_n291518# m2_26862_n291518# m2_26862_n291518# sky130_fd_pr__pfet_g5v0d10v5_CAF9E7
Xsky130_fd_pr__pfet_g5v0d10v5_CAF9E7_2 m2_27646_n292468# m2_27646_n292468# sky130_fd_sc_hvl__inv_16_1/A
+ m2_26862_n291518# m2_26862_n291518# m2_26862_n291518# sky130_fd_pr__pfet_g5v0d10v5_CAF9E7
Xsky130_fd_pr__pfet_g5v0d10v5_CAF9E7_1 m2_26866_n292108# m2_26866_n292108# m2_26960_n292468#
+ m2_26862_n291518# m2_26862_n291518# m2_26862_n291518# sky130_fd_pr__pfet_g5v0d10v5_CAF9E7
Xsky130_fd_pr__nfet_g5v0d10v5_X6E435_0 VSUBS m2_26960_n292468# m2_26960_n292468# VSUBS
+ m2_26866_n292108# m2_26866_n292108# sky130_fd_pr__nfet_g5v0d10v5_X6E435
Xsky130_fd_pr__nfet_g5v0d10v5_X6E435_2 VSUBS sky130_fd_sc_hvl__inv_16_1/A sky130_fd_sc_hvl__inv_16_1/A
+ VSUBS m2_27646_n292468# m2_27646_n292468# sky130_fd_pr__nfet_g5v0d10v5_X6E435
Xsky130_fd_pr__nfet_g5v0d10v5_X6E435_1 VSUBS m2_27646_n292468# m2_27646_n292468# VSUBS
+ m2_26960_n292468# m2_26960_n292468# sky130_fd_pr__nfet_g5v0d10v5_X6E435
Xsky130_fd_sc_hvl__inv_16_0 sky130_fd_sc_hvl__inv_16_1/A sky130_fd_sc_hvl__inv_16_0/VGND
+ VSUBS sky130_fd_sc_hvl__inv_16_1/VPB sky130_fd_sc_hvl__inv_16_0/VPWR sky130_fd_sc_hvl__inv_16_0/Y
+ sky130_fd_sc_hvl__inv_16
Xsky130_fd_sc_hvl__inv_16_1 sky130_fd_sc_hvl__inv_16_1/A sky130_fd_sc_hvl__inv_16_1/VGND
+ VSUBS sky130_fd_sc_hvl__inv_16_1/VPB sky130_fd_sc_hvl__inv_16_1/VPWR sky130_fd_sc_hvl__inv_16_1/Y
+ sky130_fd_sc_hvl__inv_16
.ends

.subckt sky130_fd_pr__pfet_01v8_X6XW7S a_63_n258# a_n33_118# a_63_118# a_n125_118#
+ a_n33_n258# a_n81_21# w_n263_n477# a_n125_n258# a_n81_n355#
X0 a_n33_n258# a_n81_n355# a_n125_n258# w_n263_n477# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X1 a_n33_118# a_n81_21# a_n125_118# w_n263_n477# sky130_fd_pr__pfet_01v8 ad=0.1155 pd=1.03 as=0.217 ps=2.02 w=0.7 l=0.15
X2 a_63_n258# a_n81_n355# a_n33_n258# w_n263_n477# sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
X3 a_63_118# a_n81_21# a_n33_118# w_n263_n477# sky130_fd_pr__pfet_01v8 ad=0.217 pd=2.02 as=0.1155 ps=1.03 w=0.7 l=0.15
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_RQPX7Z c2_n1869_n1600# m4_n1949_n1680#
X0 c2_n1869_n1600# m4_n1949_n1680# sky130_fd_pr__cap_mim_m3_2 l=16 w=16
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_HYMU45 c2_n1069_n800# m4_n1149_n880#
X0 c2_n1069_n800# m4_n1149_n880# sky130_fd_pr__cap_mim_m3_2 l=8 w=8
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_4PHTN9 m4_n1349_n1080# c2_n1269_n1000#
X0 c2_n1269_n1000# m4_n1349_n1080# sky130_fd_pr__cap_mim_m3_2 l=10 w=10
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_EEU5EF m3_n4192_n17480# c1_n4152_n17440# c1_160_n17440#
+ m3_120_n17480#
X0 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X1 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X2 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X3 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X4 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X5 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X6 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X7 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X8 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X9 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X10 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X11 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X12 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X13 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X14 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X15 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X16 c1_n4152_n17440# m3_n4192_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X17 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X18 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X19 c1_160_n17440# m3_120_n17480# sky130_fd_pr__cap_mim_m3_1 l=16 w=16
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_RRZ644 m3_n986_n840# c1_n946_n800#
X0 c1_n946_n800# m3_n986_n840# sky130_fd_pr__cap_mim_m3_1 l=8 w=8
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_KA8C77 a_516_984# a_n2292_n1416# a_n1590_n1416#
+ a_2622_984# a_1218_n1416# a_n2760_n1416# a_282_n1416# a_n654_984# a_n888_984# a_48_n1416#
+ a_n420_984# a_n420_n1416# a_750_n1416# a_n2760_984# a_1686_984# a_1452_984# a_n2526_984#
+ a_1218_984# a_n2058_n1416# a_n1356_n1416# a_2388_n1416# a_1686_n1416# a_n1824_n1416#
+ a_n2526_n1416# a_n1590_984# a_n888_n1416# a_n2890_n1546# a_516_n1416# a_n1122_984#
+ a_n1356_984# a_282_984# a_2388_984# a_2154_984# a_1920_984# a_48_984# a_n1122_n1416#
+ a_2154_n1416# a_n186_n1416# a_n186_984# a_1452_n1416# a_2622_n1416# a_1920_n1416#
+ a_984_n1416# a_n654_n1416# a_n2292_984# a_984_984# a_n1824_984# a_750_984# a_n2058_984#
X0 a_n1590_984# a_n1590_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X1 a_282_984# a_282_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X2 a_2154_984# a_2154_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X3 a_1218_984# a_1218_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X4 a_n888_984# a_n888_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X5 a_1920_984# a_1920_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X6 a_750_984# a_750_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X7 a_2622_984# a_2622_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X8 a_n2760_984# a_n2760_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X9 a_516_984# a_516_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X10 a_n186_984# a_n186_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X11 a_n2292_984# a_n2292_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X12 a_n1356_984# a_n1356_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X13 a_n2058_984# a_n2058_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X14 a_1686_984# a_1686_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X15 a_n654_984# a_n654_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X16 a_n1824_984# a_n1824_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X17 a_2388_984# a_2388_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X18 a_n420_984# a_n420_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X19 a_n2526_984# a_n2526_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X20 a_984_984# a_984_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X21 a_n1122_984# a_n1122_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X22 a_48_984# a_48_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
X23 a_1452_984# a_1452_n1416# a_n2890_n1546# sky130_fd_pr__res_xhigh_po_0p69 l=10
.ends

.subckt sky130_fd_pr__pfet_01v8_6QC8WZ a_n29_n100# a_89_n100# a_26_n197# w_n285_n319#
+ a_n92_n197# a_n147_n100#
X0 a_n29_n100# a_n92_n197# a_n147_n100# w_n285_n319# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X1 a_89_n100# a_26_n197# a_n29_n100# w_n285_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_XSEQJ6 a_189_n200# a_407_n200# a_n599_n422# a_n189_n288#
+ a_29_n288# a_247_n288# a_n407_n288# a_n29_n200# a_n247_n200# a_n465_n200#
X0 a_n247_n200# a_n407_n288# a_n465_n200# a_n599_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X1 a_407_n200# a_247_n288# a_189_n200# a_n599_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X2 a_189_n200# a_29_n288# a_n29_n200# a_n599_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X3 a_n29_n200# a_n189_n288# a_n247_n200# a_n599_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
.ends

.subckt sky130_fd_sc_ls__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=1
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0 ps=0 w=0.42 l=1
.ends

.subckt sky130_fd_sc_ls__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
X0 a_922_127# a_841_288# a_850_127# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_1598_93# a_1266_119# a_1736_119# VNB sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2 VGND a_1598_93# a_1550_119# VNB sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.0504 ps=0.66 w=0.42 l=0.15
X3 a_33_74# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.1218 ps=1.42 w=0.42 l=0.15
X4 a_1266_119# a_300_74# a_841_288# VNB sky130_fd_pr__nfet_01v8 ad=0.3067 pd=2.01 as=0.1073 ps=1.03 w=0.74 l=0.15
X5 a_1266_119# a_507_347# a_841_288# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22385 pd=1.7 as=0.39 ps=1.78 w=1 l=0.15
X6 a_714_127# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1218 pd=1.42 as=0.07245 ps=0.765 w=0.42 l=0.15
X7 a_841_288# a_714_127# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=1.78 as=0.275 ps=2.55 w=1 l=0.15
X8 VPWR a_1266_119# a_1598_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0.063 ps=0.72 w=0.42 l=0.15
X9 a_714_127# a_507_347# a_33_74# VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=0.95 as=0.1113 ps=1.37 w=0.42 l=0.15
X10 a_507_347# a_300_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.40345 pd=2.86 as=0.295 ps=2.59 w=1 l=0.15
X11 VGND RESET_B a_120_74# VNB sky130_fd_pr__nfet_01v8 ad=0.1212 pd=1.1 as=0.0504 ps=0.66 w=0.42 l=0.15
X12 VPWR a_1598_93# a_1547_508# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1550_119# a_507_347# a_1266_119# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.3067 ps=2.01 w=0.42 l=0.15
X14 a_1736_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.0819 ps=0.81 w=0.42 l=0.15
X15 a_850_127# a_300_74# a_714_127# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=0.95 w=0.42 l=0.15
X16 a_300_74# CLK_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2035 pd=2.03 as=0.1212 ps=1.1 w=0.74 l=0.15
X17 a_1547_508# a_300_74# a_1266_119# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.22385 ps=1.7 w=0.42 l=0.15
X18 a_1598_93# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0819 ps=0.81 w=0.42 l=0.15
X19 a_841_288# a_714_127# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1073 pd=1.03 as=0.24033 ps=1.715 w=0.74 l=0.15
X20 a_300_74# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.17278 ps=1.58 w=1 l=0.15
X21 VPWR a_841_288# a_817_463# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0504 ps=0.66 w=0.42 l=0.15
X22 a_120_74# D a_33_74# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X23 VPWR RESET_B a_33_74# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17278 pd=1.58 as=0.063 ps=0.72 w=0.42 l=0.15
X24 Q a_1934_94# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2146 pd=2.06 as=0.12607 ps=1.1 w=0.74 l=0.15
X25 a_817_463# a_507_347# a_714_127# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X26 VGND a_1266_119# a_1934_94# VNB sky130_fd_pr__nfet_01v8 ad=0.12607 pd=1.1 as=0.15675 ps=1.67 w=0.55 l=0.15
X27 a_714_127# a_300_74# a_33_74# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X28 VGND RESET_B a_922_127# VNB sky130_fd_pr__nfet_01v8 ad=0.24033 pd=1.715 as=0.0441 ps=0.63 w=0.42 l=0.15
X29 a_507_347# a_300_74# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2479 pd=2.15 as=0.3299 ps=2.67 w=0.74 l=0.15
X30 VPWR a_1266_119# a_1934_94# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1862 pd=1.475 as=0.231 ps=2.23 w=0.84 l=0.15
X31 Q a_1934_94# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3192 pd=2.81 as=0.1862 ps=1.475 w=1.12 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_XJT6XQ a_n33_n50# a_63_n50# a_n125_n50# a_n81_n157#
+ w_n263_n269#
X0 a_n33_n50# a_n81_n157# a_n125_n50# w_n263_n269# sky130_fd_pr__pfet_01v8 ad=0.0825 pd=0.83 as=0.155 ps=1.62 w=0.5 l=0.15
X1 a_63_n50# a_n81_n157# a_n33_n50# w_n263_n269# sky130_fd_pr__pfet_01v8 ad=0.155 pd=1.62 as=0.0825 ps=0.83 w=0.5 l=0.15
.ends

.subckt TieH_1p8 TieH VSS VCC
XXM4 VSS m2_456_n646# m2_456_n646# VSS sky130_fd_pr__nfet_01v8_L9ESAD
XXM5 TieH VCC VCC m2_456_n646# VCC sky130_fd_pr__pfet_01v8_XJT6XQ
.ends

.subckt sky130_fd_sc_ls__buf_8 A VGND VNB VPB VPWR X
X0 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8 ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8 ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5 VPWR A a_27_74# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X7 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8 ad=0.12025 pd=1.065 as=0.2109 ps=2.05 w=0.74 l=0.15
X8 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8 ad=0.2627 pd=2.19 as=0.10545 ps=1.025 w=0.74 l=0.15
X9 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X10 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.12025 ps=1.065 w=0.74 l=0.15
X11 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3304 pd=2.83 as=0.1764 ps=1.435 w=1.12 l=0.15
X12 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8 ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X13 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X14 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1876 pd=1.455 as=0.168 ps=1.42 w=1.12 l=0.15
X15 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10545 pd=1.025 as=0.1554 ps=1.16 w=0.74 l=0.15
X16 VPWR A a_27_74# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X17 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X18 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X19 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X20 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X21 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.435 as=0.1876 ps=1.455 w=1.12 l=0.15
.ends

.subckt sky130_fd_sc_ls__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 VPWR RESET_B a_30_78# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.05985 ps=0.705 w=0.42 l=0.15
X1 VGND RESET_B a_894_138# VNB sky130_fd_pr__nfet_01v8 ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2 a_894_138# a_830_359# a_816_138# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X3 VPWR a_1518_203# a_1468_493# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_1864_409# a_1266_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X5 a_830_359# a_695_457# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X6 a_816_138# a_490_390# a_695_457# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X7 a_1476_81# a_306_96# a_1266_74# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X8 VGND a_1864_409# Q VNB sky130_fd_pr__nfet_01v8 ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X9 a_490_390# a_306_96# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.15 ps=1.3 w=1 l=0.15
X10 a_1468_493# a_490_390# a_1266_74# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X11 VPWR CLK a_306_96# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.31 ps=2.62 w=1 l=0.15
X12 a_1266_74# a_306_96# a_830_359# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X13 a_830_359# a_695_457# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X14 VPWR a_1864_409# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X15 a_1656_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X16 VPWR a_1266_74# a_1518_203# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X17 a_1864_409# a_1266_74# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X18 VGND CLK a_306_96# VNB sky130_fd_pr__nfet_01v8 ad=0.16238 pd=1.255 as=0.2646 ps=2.4 w=0.74 l=0.15
X19 a_1518_203# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X20 a_695_457# a_306_96# a_30_78# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X21 a_1518_203# a_1266_74# a_1656_81# VNB sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X22 a_695_457# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X23 a_117_78# D a_30_78# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X24 VPWR a_830_359# a_785_457# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X25 VGND a_1518_203# a_1476_81# VNB sky130_fd_pr__nfet_01v8 ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X26 VGND RESET_B a_117_78# VNB sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X27 a_785_457# a_306_96# a_695_457# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X28 a_695_457# a_490_390# a_30_78# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.1218 ps=1.42 w=0.42 l=0.15
X29 a_30_78# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05985 pd=0.705 as=0.1197 ps=1.41 w=0.42 l=0.15
X30 a_490_390# a_306_96# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2183 pd=2.07 as=0.16238 ps=1.255 w=0.74 l=0.15
X31 a_1266_74# a_490_390# a_830_359# VNB sky130_fd_pr__nfet_01v8 ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
.ends

.subckt sky130_fd_sc_ls__xor2_1 A B VGND VNB VPB VPWR X
X0 X B a_455_87# VNB sky130_fd_pr__nfet_01v8 ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X1 X a_194_125# a_355_368# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
X2 a_194_125# B a_158_392# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A a_355_368# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2352 pd=1.54 as=0.3752 ps=2.91 w=1.12 l=0.15
X4 a_158_392# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X5 a_355_368# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.196 pd=1.47 as=0.2352 ps=1.54 w=1.12 l=0.15
X6 a_194_125# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17738 pd=1.195 as=0.33275 ps=2.31 w=0.55 l=0.15
X7 a_455_87# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0888 pd=0.98 as=0.12607 ps=1.1 w=0.74 l=0.15
X8 VGND B a_194_125# VNB sky130_fd_pr__nfet_01v8 ad=0.12607 pd=1.1 as=0.17738 ps=1.195 w=0.55 l=0.15
X9 VGND a_194_125# X VNB sky130_fd_pr__nfet_01v8 ad=0.2997 pd=2.29 as=0.1554 ps=1.16 w=0.74 l=0.15
.ends

.subckt delayPulse_digital sky130_fd_sc_ls__dfrtp_1_0/RESET_B sky130_fd_sc_ls__dfrtp_1_0/CLK
+ sky130_fd_sc_ls__dfrtn_1_0/Q sky130_fd_sc_ls__dfrtp_1_0/Q sky130_fd_sc_ls__xor2_1_0/B
+ sky130_fd_sc_ls__xor2_1_0/A TieH_1p8_0/VCC VSUBS
Xsky130_fd_sc_ls__decap_4_0 VSUBS VSUBS TieH_1p8_0/VCC TieH_1p8_0/VCC sky130_fd_sc_ls__decap_4
Xsky130_fd_sc_ls__dfrtn_1_0 sky130_fd_sc_ls__buf_8_0/X TieH_1p8_0/TieH sky130_fd_sc_ls__dfrtp_1_0/CLK
+ VSUBS VSUBS TieH_1p8_0/VCC TieH_1p8_0/VCC sky130_fd_sc_ls__dfrtn_1_0/Q sky130_fd_sc_ls__dfrtn_1
XTieH_1p8_0 TieH_1p8_0/TieH VSUBS TieH_1p8_0/VCC TieH_1p8
Xsky130_fd_sc_ls__buf_8_0 sky130_fd_sc_ls__buf_8_0/A VSUBS VSUBS TieH_1p8_0/VCC TieH_1p8_0/VCC
+ sky130_fd_sc_ls__buf_8_0/X sky130_fd_sc_ls__buf_8
Xsky130_fd_sc_ls__dfrtp_1_0 sky130_fd_sc_ls__dfrtp_1_0/CLK TieH_1p8_0/TieH sky130_fd_sc_ls__dfrtp_1_0/RESET_B
+ VSUBS VSUBS TieH_1p8_0/VCC TieH_1p8_0/VCC sky130_fd_sc_ls__dfrtp_1_0/Q sky130_fd_sc_ls__dfrtp_1
Xsky130_fd_sc_ls__xor2_1_0 sky130_fd_sc_ls__xor2_1_0/A sky130_fd_sc_ls__xor2_1_0/B
+ VSUBS VSUBS TieH_1p8_0/VCC TieH_1p8_0/VCC sky130_fd_sc_ls__buf_8_0/A sky130_fd_sc_ls__xor2_1
.ends

.subckt delayPulse_final din por porb porb_h[0] porb_h[1] ibn180n m2_1725_n286520#
+ VCCH VCCL m2_1729_n290386# VSS VT2
XXM12 VT3 VCCL VT2 VCCL VT2 VCCL sky130_fd_pr__pfet_01v8_GHZ9W9
XXM23 m2_27024_n287466# m2_27024_n287466# vbp1 vbp1 m2_27024_n287466# VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXM34 VSS VSS m4_25183_n288425# m2_24504_n284758# sky130_fd_pr__nfet_01v8_L9ESAD
Xsky130_fd_pr__cap_mim_m3_2_2V27AY_0 VT3 VCCL VCCL VT3 sky130_fd_pr__cap_mim_m3_2_2V27AY
Xpor_output_buffer_1 VCCL por VSS porPre por_output_buffer
XXM13 m2_31224_n287586# VT3 VSS VSS VSS VT3 sky130_fd_pr__nfet_01v8_G7LLWL
XXM24 ibn180n ibn180n VCCH m1_22999_n287228# sky130_fd_pr__pfet_g5v0d10v5_PQJ659
XXM35 VCCL m4_25183_n288425# VCCL VCCL m2_24504_n284758# m4_25183_n288425# m2_24504_n284758#
+ sky130_fd_pr__pfet_01v8_U6B66J
Xsky130_fd_pr__cap_mim_m3_2_2V27AY_1 VT2 VSS VSS VT2 sky130_fd_pr__cap_mim_m3_2_2V27AY
XXM14 m2_27024_n287466# m2_31224_n287586# VT3 VT3 m2_27024_n287466# m2_31224_n287586#
+ m2_27024_n287466# sky130_fd_pr__pfet_01v8_SKYQWJ
XXM25 m1_22999_n287228# m1_22999_n287228# m1_22999_n287228# m1_22999_n287228# VCCH
+ m1_22999_n287228# m1_22999_n287228# m1_22999_n287228# VCCH m1_22999_n287228# m1_22999_n287228#
+ m1_22999_n287228# m1_22999_n287228# VCCH VCCH VCCH m1_22999_n287228# VCCH sky130_fd_pr__pfet_g5v0d10v5_KLZS5A
XXM36 VSS VSS Td_Sd Td_Sd m2_24748_n284671# sky130_fd_pr__nfet_01v8_5QNSAB
Xx3 porbPre x3/aout VCCL VSS VCCH levelShifter
XXM26 m1_22125_n286949# VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5_69TNYL
XXM16 m2_27024_n287466# VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXM27 VSS VSS m2_31224_n287586# m2_31884_n287663# sky130_fd_pr__nfet_01v8_L9ESAD
XXM38 VSS VSS m2_24504_n284758# m2_24748_n284671# sky130_fd_pr__nfet_01v8_L9ESAD
XXM17 VSS vbp1 VSS vbn1 sky130_fd_pr__nfet_g5v0d10v5_ESEQJ8
XXM39 VCCL m2_24504_n284758# VCCL VCCL m2_24748_n284671# m2_24504_n284758# m2_24748_n284671#
+ sky130_fd_pr__pfet_01v8_U6B66J
Xsky130_fd_pr__cap_mim_m3_1_TBT74C_0 vbp1 VCCL sky130_fd_pr__cap_mim_m3_1_TBT74C
XXM18 m1_22999_n287228# VCCH VCCH m2_24152_n287606# sky130_fd_pr__pfet_g5v0d10v5_PQJ659
XXM29 VCCL m2_31224_n287586# VCCL VCCL m2_31884_n287663# m2_31224_n287586# m2_31884_n287663#
+ sky130_fd_pr__pfet_01v8_U6B66J
Xsky130_fd_pr__cap_mim_m3_1_TBT74C_1 vbn1 VSS sky130_fd_pr__cap_mim_m3_1_TBT74C
XXM19 vbn1 VSS vbn1 VSS VSS vbn1 vbn1 vbn1 vbn1 vbn1 vbn1 vbn1 VSS vbn1 VSS vbn1 sky130_fd_pr__nfet_g5v0d10v5_SYBQJL
Xsky130_fd_pr__cap_mim_m3_1_TBT74C_2 m1_22999_n287228# VCCH sky130_fd_pr__cap_mim_m3_1_TBT74C
XXM1 vbp1 VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
Xsky130_fd_pr__cap_mim_m3_1_KB5CJD_0 VCCL m4_25183_n288425# sky130_fd_pr__cap_mim_m3_1_KB5CJD
XXM2 VCCL m2_30306_n287752# din din VCCL m2_30306_n287752# VCCL sky130_fd_pr__pfet_01v8_SKYQWJ
Xsky130_fd_pr__cap_mim_m3_1_KB5CJD_1 VCCL m2_24748_n284671# sky130_fd_pr__cap_mim_m3_1_KB5CJD
XXM3 VCCL Td_S m2_30306_n287752# m2_30306_n287752# VCCL Td_S VCCL sky130_fd_pr__pfet_01v8_SKYQWJ
Xsky130_fd_pr__cap_mim_m3_1_KB5CJD_2 VSS m2_24504_n284758# sky130_fd_pr__cap_mim_m3_1_KB5CJD
XXM4 Td_Lb VSS VSS VSS Td_L sky130_fd_pr__nfet_01v8_5QNSAB
XXM5 VT2 m2_30306_n287752# VSS VSS VSS m2_30306_n287752# sky130_fd_pr__nfet_01v8_G7LLWL
XXM6 VT3 VT2 VSS m2_29342_n288187# m2_29342_n288187# VT2 sky130_fd_pr__nfet_01v8_G7LLWL
Xpor_output_driver_h_0 VCCH porb_h[0] VCCH VSS VCCH x3/aout VCCH VSS porb_h[1] VSS
+ por_output_driver_h
XXM7 VSS din VSS m2_30306_n287752# m2_30306_n287752# din sky130_fd_pr__nfet_01v8_G7LLWL
XXM8 VSS m2_30306_n287752# VSS Td_S Td_S m2_30306_n287752# sky130_fd_pr__nfet_01v8_G7LLWL
XXM9 VCCL Td_Lb VCCL VCCL Td_Lb Td_L VCCL VCCL Td_L sky130_fd_pr__pfet_01v8_X6XW7S
Xsky130_fd_pr__cap_mim_m3_2_RQPX7Z_0 VCCL vbp1 sky130_fd_pr__cap_mim_m3_2_RQPX7Z
XXC1 VSS vbn1 sky130_fd_pr__cap_mim_m3_2_RQPX7Z
Xsky130_fd_pr__pfet_01v8_XPC8Y6_1[0] vbp1 VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
Xsky130_fd_pr__pfet_01v8_XPC8Y6_1[1] vbp1 VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
Xsky130_fd_pr__pfet_01v8_XPC8Y6_1[2] vbp1 VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
Xsky130_fd_pr__pfet_01v8_XPC8Y6_1[3] vbp1 VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
Xsky130_fd_pr__pfet_01v8_XPC8Y6_1[4] vbp1 VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
Xsky130_fd_pr__pfet_01v8_XPC8Y6_1[5] VCCL m2_29064_n286804# vbp1 vbp1 m2_29064_n286804#
+ VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
Xsky130_fd_pr__pfet_01v8_XPC8Y6_1[6] m2_29064_n286804# m2_29064_n286804# vbp1 vbp1
+ m2_29064_n286804# VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXC3 VCCH ibn180n sky130_fd_pr__cap_mim_m3_2_HYMU45
XXC4 m4_25183_n288425# VCCL sky130_fd_pr__cap_mim_m3_2_4PHTN9
XXC5 VCCH m1_22999_n287228# sky130_fd_pr__cap_mim_m3_2_RQPX7Z
Xsky130_fd_pr__cap_mim_m3_2_4PHTN9_0 m2_24504_n284758# VSS sky130_fd_pr__cap_mim_m3_2_4PHTN9
Xsky130_fd_pr__cap_mim_m3_1_EEU5EF_0 VSS VT2 VT2 VSS sky130_fd_pr__cap_mim_m3_1_EEU5EF
XXC9 m2_24748_n284671# VCCL sky130_fd_pr__cap_mim_m3_2_4PHTN9
Xsky130_fd_pr__cap_mim_m3_1_EEU5EF_1 VCCL VT3 VT3 VCCL sky130_fd_pr__cap_mim_m3_1_EEU5EF
Xsky130_fd_pr__cap_mim_m3_1_RRZ644_0 VCCH ibn180n sky130_fd_pr__cap_mim_m3_1_RRZ644
XXM40 Td_Sd VCCL Td_Sd Td_Sd VCCL m2_24748_n284671# VCCL Td_Sd m2_24748_n284671# sky130_fd_pr__pfet_01v8_X6XW7S
XXM30 Td_L VSS VSS VSS m2_31884_n287663# sky130_fd_pr__nfet_01v8_5QNSAB
XXM20 vbp1 VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXM31 VCCL Td_L VCCL VCCL Td_L m2_31884_n287663# VCCL VCCL m2_31884_n287663# sky130_fd_pr__pfet_01v8_X6XW7S
Xsky130_fd_pr__res_xhigh_po_0p69_KA8C77_2 m1_19785_n286949# m1_17211_n289349# m1_17679_n289349#
+ m1_22125_n286949# m1_20487_n289349# m1_16743_n289349# m1_19551_n289349# m1_18849_n286949#
+ m1_18381_n286949# m1_19551_n289349# m1_18849_n286949# m1_19083_n289349# m1_20019_n289349#
+ m1_16739_n286950# m1_21189_n286949# m1_20721_n286949# m1_16977_n286949# m1_20721_n286949#
+ m1_17211_n289349# m1_18147_n289349# m1_21891_n289349# m1_20955_n289349# m1_17679_n289349#
+ m1_16743_n289349# m1_17913_n286949# m1_18615_n289349# VSS m1_20019_n289349# m1_18381_n286949#
+ m1_17913_n286949# m1_19785_n286949# m1_21657_n286949# m1_21657_n286949# m1_21189_n286949#
+ m1_19317_n286949# m1_18147_n289349# m1_21423_n289349# m1_19083_n289349# m1_19317_n286949#
+ m1_20955_n289349# m1_21891_n289349# m1_21423_n289349# m1_20487_n289349# m1_18615_n289349#
+ m1_16977_n286949# m1_20253_n286949# m1_17445_n286949# m1_20253_n286949# m1_17445_n286949#
+ sky130_fd_pr__res_xhigh_po_0p69_KA8C77
XXM10 VT2 m2_29064_n286804# m2_30306_n287752# VCCL m2_30306_n287752# m2_29064_n286804#
+ sky130_fd_pr__pfet_01v8_6QC8WZ
XXM21 VSS m2_29342_n288187# VSS vbn1 vbn1 vbn1 vbn1 m2_29342_n288187# VSS m2_29342_n288187#
+ sky130_fd_pr__nfet_g5v0d10v5_XSEQJ6
XXM32 VSS VSS Td_S m4_25183_n288425# sky130_fd_pr__nfet_01v8_L9ESAD
XdelayPulse_digital_0 Td_Lb Td_Sd porbPre porPre Td_Sd Td_L VCCL VSS delayPulse_digital
Xsky130_fd_pr__res_xhigh_po_0p69_KA8C77_3 m1_20018_n283415# m1_16975_n285816# m1_17911_n285816#
+ m1_21890_n283415# m1_20719_n285816# m1_16739_n286950# m1_19783_n285816# m1_18614_n283415#
+ m1_18614_n283415# m1_19315_n285816# m1_19082_n283415# m1_18847_n285816# m1_20251_n285816#
+ m1_16742_n283415# m1_20954_n283415# m1_20954_n283415# m1_16742_n283415# m1_20486_n283415#
+ m1_17443_n285816# m1_17911_n285816# m1_21655_n285816# m1_21187_n285816# m1_17443_n285816#
+ m1_16975_n285816# m1_17678_n283415# m1_18379_n285816# VSS m1_19783_n285816# m1_18146_n283415#
+ m1_18146_n283415# m1_19550_n283415# m1_21890_n283415# m1_21422_n283415# m1_21422_n283415#
+ m1_19550_n283415# m1_18379_n285816# m1_21655_n285816# m1_19315_n285816# m1_19082_n283415#
+ m1_20719_n285816# VSS m1_21187_n285816# m1_20251_n285816# m1_18847_n285816# m1_17210_n283415#
+ m1_20486_n283415# m1_17678_n283415# m1_20018_n283415# m1_17210_n283415# sky130_fd_pr__res_xhigh_po_0p69_KA8C77
XXM11 ibn180n m2_24152_n287606# VCCH vbn1 sky130_fd_pr__pfet_g5v0d10v5_PQJ659
XXM22[0] m2_27024_n287466# VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXM22[1] m2_27024_n287466# VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXM22[2] m2_27024_n287466# VCCL vbp1 vbp1 VCCL VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXM22[3] vbp1 vbp1 vbp1 vbp1 vbp1 VCCL sky130_fd_pr__pfet_01v8_XPC8Y6
XXM33 VCCL Td_S VCCL VCCL m4_25183_n288425# Td_S m4_25183_n288425# sky130_fd_pr__pfet_01v8_U6B66J
Xpor_output_buffer_0 VCCL porb VSS porbPre por_output_buffer
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_WGPHGK a_1625_n4416# a_463_3984# a_n699_3984#
+ a_n2157_n4546# a_n1197_3984# a_n1363_n4416# a_297_3984# a_1127_n4416# a_n533_n4416#
+ a_1957_3984# a_n1861_3984# a_961_3984# a_n35_n4416# a_795_n4416# a_n1695_3984# a_1957_n4416#
+ a_795_3984# a_n201_3984# a_n1695_n4416# a_n2027_3984# a_n1529_3984# a_297_n4416#
+ a_1459_n4416# a_629_3984# a_n35_3984# a_n865_n4416# a_629_n4416# a_1293_3984# a_n1197_n4416#
+ a_n367_n4416# a_n1529_n4416# a_n533_3984# a_131_n4416# a_n1031_3984# a_1127_3984#
+ a_n2027_n4416# a_131_3984# a_n367_3984# a_1791_3984# a_n1031_n4416# a_1791_n4416#
+ a_961_n4416# a_n201_n4416# a_1625_3984# a_n699_n4416# a_n865_3984# a_n1861_n4416#
+ a_1459_3984# a_1293_n4416# a_463_n4416# a_n1363_3984#
X0 a_n1197_3984# a_n1197_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X1 a_n1695_3984# a_n1695_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X2 a_n533_3984# a_n533_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X3 a_1127_3984# a_1127_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X4 a_463_3984# a_463_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X5 a_629_3984# a_629_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X6 a_n1031_3984# a_n1031_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X7 a_n35_3984# a_n35_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X8 a_1625_3984# a_1625_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X9 a_961_3984# a_961_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X10 a_n367_3984# a_n367_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X11 a_297_3984# a_297_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X12 a_n865_3984# a_n865_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X13 a_1293_3984# a_1293_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X14 a_1459_3984# a_1459_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X15 a_795_3984# a_795_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X16 a_n1529_3984# a_n1529_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X17 a_n2027_3984# a_n2027_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X18 a_n1363_3984# a_n1363_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X19 a_1791_3984# a_1791_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X20 a_1957_3984# a_1957_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X21 a_n201_3984# a_n201_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X22 a_n1861_3984# a_n1861_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X23 a_n699_3984# a_n699_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X24 a_131_3984# a_131_n4416# a_n2157_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_FPTPS4 a_n90_n188# a_90_n100# a_n282_n322# a_n148_n100#
X0 a_90_n100# a_n90_n188# a_n148_n100# a_n282_n322# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.9
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_CZFQWY a_90_n309# a_n90_21# a_n148_n309# a_n282_n531#
+ a_n148_109# a_90_109# a_n90_n397#
X0 a_90_109# a_n90_21# a_n148_109# a_n282_n531# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.9
X1 a_90_n309# a_n90_n397# a_n148_n309# a_n282_n531# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.9
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_PXB2PH a_214_n4016# a_n284_3584# a_48_n4016#
+ a_n118_3584# a_n284_n4016# a_214_3584# a_n414_n4146# a_n118_n4016# a_48_3584#
X0 a_n284_3584# a_n284_n4016# a_n414_n4146# sky130_fd_pr__res_xhigh_po_0p35 l=36
X1 a_48_3584# a_48_n4016# a_n414_n4146# sky130_fd_pr__res_xhigh_po_0p35 l=36
X2 a_214_3584# a_214_n4016# a_n414_n4146# sky130_fd_pr__res_xhigh_po_0p35 l=36
X3 a_n118_3584# a_n118_n4016# a_n414_n4146# sky130_fd_pr__res_xhigh_po_0p35 l=36
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_MNWQZD a_463_3984# a_n699_3984# a_n1197_3984#
+ a_297_3984# a_1127_n4416# a_n533_n4416# a_961_3984# a_n35_n4416# a_795_n4416# a_795_3984#
+ a_n201_3984# a_297_n4416# a_629_3984# a_n35_3984# a_n865_n4416# a_629_n4416# a_n1197_n4416#
+ a_n367_n4416# a_n533_3984# a_n1327_n4546# a_131_n4416# a_n1031_3984# a_1127_3984#
+ a_131_3984# a_n367_3984# a_n1031_n4416# a_961_n4416# a_n201_n4416# a_n699_n4416#
+ a_n865_3984# a_463_n4416#
X0 a_n1197_3984# a_n1197_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X1 a_n533_3984# a_n533_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X2 a_1127_3984# a_1127_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X3 a_463_3984# a_463_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X4 a_629_3984# a_629_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X5 a_n1031_3984# a_n1031_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X6 a_n35_3984# a_n35_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X7 a_961_3984# a_961_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X8 a_n367_3984# a_n367_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X9 a_297_3984# a_297_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X10 a_n865_3984# a_n865_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X11 a_795_3984# a_795_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X12 a_n201_3984# a_n201_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X13 a_n699_3984# a_n699_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
X14 a_131_3984# a_131_n4416# a_n1327_n4546# sky130_fd_pr__res_xhigh_po_0p35 l=40
.ends

.subckt sky130_sw_ip__por por avdd dvdd porb dvss porb_h[0] porb_h[1] avss
Xx1 x1/Vinn x1/Vinp x2/din avdd dvdd x2/ibn180n x1/vo avss comparator_final
Xx2 x2/din por porb porb_h[0] porb_h[1] x2/ibn180n avdd avdd dvdd avss dvss x2/VT2
+ delayPulse_final
XR1 m1_10763_n288829# m1_9601_n280429# m1_8273_n280429# avss m1_7941_n280429# m1_7775_n288829#
+ m1_9269_n280429# m1_10099_n288829# m1_8439_n288829# m1_10929_n280429# m1_7277_n280429#
+ m1_9933_n280429# m1_9103_n288829# m1_9767_n288829# m1_7277_n280429# x1/Vinn m1_9933_n280429#
+ m1_8937_n280429# m1_7443_n288829# avss m1_7609_n280429# m1_9435_n288829# m1_10431_n288829#
+ m1_9601_n280429# m1_8937_n280429# m1_8107_n288829# m1_9767_n288829# m1_10265_n280429#
+ m1_7775_n288829# m1_8771_n288829# m1_7443_n288829# m1_8605_n280429# m1_9103_n288829#
+ m1_7941_n280429# m1_10265_n280429# m1_7111_n288829# m1_9269_n280429# m1_8605_n280429#
+ m1_10929_n280429# m1_8107_n288829# m1_10763_n288829# m1_10099_n288829# m1_8771_n288829#
+ m1_10597_n280429# m1_8439_n288829# m1_8273_n280429# m1_7111_n288829# m1_10597_n280429#
+ m1_10431_n288829# m1_9435_n288829# m1_7609_n280429# sky130_fd_pr__res_xhigh_po_0p35_WGPHGK
Xsky130_fd_pr__nfet_05v0_nvt_FPTPS4_0 x1/vo m2_10326_n290222# avss x1/Vinn sky130_fd_pr__nfet_05v0_nvt_FPTPS4
XXM2 m1_15791_n280880# avdd avdd avss m1_14983_n280431# m1_15791_n280880# avdd sky130_fd_pr__nfet_05v0_nvt_CZFQWY
XR10 x1/Vinp m1_11633_n281148# m2_10326_n290222# m1_11633_n281148# x1/Vinn m1_11964_n281149#
+ avss x1/Vinp m1_11964_n281149# sky130_fd_pr__res_xhigh_po_0p35_PXB2PH
XR12 m1_14304_n280429# m1_12968_n280429# m1_12634_n280429# m1_13970_n280429# m1_14804_n288829#
+ m1_13134_n288829# m1_14638_n280429# m1_13802_n288829# m1_14470_n288829# m1_14638_n280429#
+ m1_13636_n280429# m1_14136_n288829# m1_14304_n280429# m1_13636_n280429# m1_12800_n288829#
+ m1_14470_n288829# x1/Vinp m1_13468_n288829# m1_13302_n280429# avss m1_13802_n288829#
+ m1_12634_n280429# m1_14983_n280431# m1_13970_n280429# m1_13302_n280429# m1_12800_n288829#
+ m1_14804_n288829# m1_13468_n288829# m1_13134_n288829# m1_12968_n280429# m1_14136_n288829#
+ sky130_fd_pr__res_xhigh_po_0p35_MNWQZD
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_SABQJA a_n345_n200# a_129_n200# a_n503_n200#
+ a_287_n200# a_445_n200# a_n637_n422# a_29_n288# a_n129_n288# a_187_n288# a_n287_n288#
+ a_345_n288# a_n29_n200# a_n187_n200# a_n445_n288#
X0 a_n187_n200# a_n287_n288# a_n345_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X1 a_287_n200# a_187_n288# a_129_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X2 a_n345_n200# a_n445_n288# a_n503_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X3 a_129_n200# a_29_n288# a_n29_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X4 a_445_n200# a_345_n288# a_287_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X5 a_n29_n200# a_n129_n288# a_n187_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_LQS9ZD a_n819_n200# a_n345_n200# a_n977_n200#
+ a_29_n297# a_n129_n297# a_187_n297# a_129_n200# a_n503_n200# a_n287_n297# a_819_n297#
+ a_345_n297# a_287_n200# a_n661_n200# a_n919_n297# w_n1177_n497# a_n445_n297# a_919_n200#
+ a_503_n297# a_445_n200# a_n603_n297# a_661_n297# a_603_n200# a_n761_n297# a_761_n200#
+ a_n29_n200# a_n187_n200#
X0 a_n819_n200# a_n919_n297# a_n977_n200# w_n1177_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X1 a_n661_n200# a_n761_n297# a_n819_n200# w_n1177_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X2 a_919_n200# a_819_n297# a_761_n200# w_n1177_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X3 a_n187_n200# a_n287_n297# a_n345_n200# w_n1177_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X4 a_761_n200# a_661_n297# a_603_n200# w_n1177_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X5 a_287_n200# a_187_n297# a_129_n200# w_n1177_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X6 a_n345_n200# a_n445_n297# a_n503_n200# w_n1177_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X7 a_129_n200# a_29_n297# a_n29_n200# w_n1177_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X8 a_445_n200# a_345_n297# a_287_n200# w_n1177_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X9 a_n503_n200# a_n603_n297# a_n661_n200# w_n1177_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X10 a_n29_n200# a_n129_n297# a_n187_n200# w_n1177_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X11 a_603_n200# a_503_n297# a_445_n200# w_n1177_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EJGQJV a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt isolated_switch_3 on off vdd shunt vss out in
XXM15 m2_961_43# in in m2_961_43# in vss on on on on on m2_961_43# in on sky130_fd_pr__nfet_g5v0d10v5_SABQJA
Xsky130_fd_pr__pfet_g5v0d10v5_LQS9ZD_0 m2_961_43# out out off off off m2_961_43# m2_961_43#
+ off off off out out off vdd off out off m2_961_43# off off out off m2_961_43# out
+ m2_961_43# sky130_fd_pr__pfet_g5v0d10v5_LQS9ZD
XXM4 in m2_961_43# m2_961_43# off off off in in off off off m2_961_43# m2_961_43#
+ off vdd off m2_961_43# off in off off m2_961_43# off in m2_961_43# in sky130_fd_pr__pfet_g5v0d10v5_LQS9ZD
Xsky130_fd_pr__nfet_g5v0d10v5_SABQJA_0 out m2_961_43# m2_961_43# out m2_961_43# vss
+ on on on on on out m2_961_43# on sky130_fd_pr__nfet_g5v0d10v5_SABQJA
Xsky130_fd_pr__nfet_g5v0d10v5_EJGQJV_0 vss vss m2_961_43# shunt sky130_fd_pr__nfet_g5v0d10v5_EJGQJV
.ends

.subckt isolated_switch_large avss on avdd off dvdd out in dvss
Xx2 on dvdd dvss avdd avdd x2/X avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xx3 off dvdd dvss avdd avdd x3/X avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__diode_2_0 off dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xisolated_switch_3_0 x2/X isolated_switch_3_0/off avdd x3/X avss out in isolated_switch_3
Xsky130_fd_sc_hvl__diode_2_1 on dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_1_0 x2/X dvss dvss avdd avdd isolated_switch_3_0/off sky130_fd_sc_hvl__inv_1
.ends

.subckt switch_array_18 isolated_switch_large_0[1|0]/on right_instramp_out isolated_switch_large_0[1|2]/off
+ left_instramp_out isolated_switch_large_0[5|1]/on isolated_switch_large_0[5|0]/on
+ right_hgbw_opamp_out isolated_switch_large_0[2|2]/on isolated_switch_large_0[2|1]/off
+ dvdd dvss isolated_switch_large_0[4|0]/off isolated_switch_large_0[4|2]/on isolated_switch_large_0[0|0]/on
+ avdd isolated_switch_large_0[1|0]/off isolated_switch_large_0[5|2]/on isolated_switch_large_0[5|0]/off
+ isolated_switch_large_0[3|1]/off isolated_switch_large_0[3|2]/on left_hgbw_opamp_out
+ isolated_switch_large_0[3|1]/on isolated_switch_large_0[0|1]/off isolated_switch_large_0[0|1]/on
+ comp_p isolated_switch_large_0[2|1]/on adc0 isolated_switch_large_0[0|0]/off isolated_switch_large_0[1|1]/off
+ isolated_switch_large_0[4|0]/on isolated_switch_large_0[4|1]/on isolated_switch_large_0[4|1]/off
+ isolated_switch_large_0[2|0]/off isolated_switch_large_0[3|0]/on isolated_switch_large_0[5|1]/off
+ comp_n isolated_switch_large_0[3|2]/off ulpcomp_p isolated_switch_large_0[0|2]/off
+ adc1 isolated_switch_large_0[3|0]/off isolated_switch_large_0[5|2]/off ulpcomp_n
+ isolated_switch_large_0[2|0]/on right_lp_opamp_out isolated_switch_large_0[2|2]/off
+ isolated_switch_large_0[1|1]/on isolated_switch_large_0[4|2]/off isolated_switch_large_0[1|2]/on
+ left_lp_opamp_out isolated_switch_large_0[0|2]/on avss
Xisolated_switch_large_0[0|0] avss isolated_switch_large_0[0|0]/on avdd isolated_switch_large_0[0|0]/off
+ dvdd left_lp_opamp_out ulpcomp_n dvss isolated_switch_large
Xisolated_switch_large_0[1|0] avss isolated_switch_large_0[1|0]/on avdd isolated_switch_large_0[1|0]/off
+ dvdd left_lp_opamp_out comp_n dvss isolated_switch_large
Xisolated_switch_large_0[2|0] avss isolated_switch_large_0[2|0]/on avdd isolated_switch_large_0[2|0]/off
+ dvdd left_lp_opamp_out adc1 dvss isolated_switch_large
Xisolated_switch_large_0[3|0] avss isolated_switch_large_0[3|0]/on avdd isolated_switch_large_0[3|0]/off
+ dvdd right_lp_opamp_out ulpcomp_p dvss isolated_switch_large
Xisolated_switch_large_0[4|0] avss isolated_switch_large_0[4|0]/on avdd isolated_switch_large_0[4|0]/off
+ dvdd right_lp_opamp_out comp_p dvss isolated_switch_large
Xisolated_switch_large_0[5|0] avss isolated_switch_large_0[5|0]/on avdd isolated_switch_large_0[5|0]/off
+ dvdd right_lp_opamp_out adc0 dvss isolated_switch_large
Xisolated_switch_large_0[0|1] avss isolated_switch_large_0[0|1]/on avdd isolated_switch_large_0[0|1]/off
+ dvdd right_hgbw_opamp_out ulpcomp_n dvss isolated_switch_large
Xisolated_switch_large_0[1|1] avss isolated_switch_large_0[1|1]/on avdd isolated_switch_large_0[1|1]/off
+ dvdd right_hgbw_opamp_out comp_n dvss isolated_switch_large
Xisolated_switch_large_0[2|1] avss isolated_switch_large_0[2|1]/on avdd isolated_switch_large_0[2|1]/off
+ dvdd right_hgbw_opamp_out adc1 dvss isolated_switch_large
Xisolated_switch_large_0[3|1] avss isolated_switch_large_0[3|1]/on avdd isolated_switch_large_0[3|1]/off
+ dvdd left_hgbw_opamp_out ulpcomp_p dvss isolated_switch_large
Xisolated_switch_large_0[4|1] avss isolated_switch_large_0[4|1]/on avdd isolated_switch_large_0[4|1]/off
+ dvdd left_hgbw_opamp_out comp_p dvss isolated_switch_large
Xisolated_switch_large_0[5|1] avss isolated_switch_large_0[5|1]/on avdd isolated_switch_large_0[5|1]/off
+ dvdd left_hgbw_opamp_out adc0 dvss isolated_switch_large
Xisolated_switch_large_0[0|2] avss isolated_switch_large_0[0|2]/on avdd isolated_switch_large_0[0|2]/off
+ dvdd right_instramp_out ulpcomp_n dvss isolated_switch_large
Xisolated_switch_large_0[1|2] avss isolated_switch_large_0[1|2]/on avdd isolated_switch_large_0[1|2]/off
+ dvdd right_instramp_out comp_n dvss isolated_switch_large
Xisolated_switch_large_0[2|2] avss isolated_switch_large_0[2|2]/on avdd isolated_switch_large_0[2|2]/off
+ dvdd right_instramp_out adc1 dvss isolated_switch_large
Xisolated_switch_large_0[3|2] avss isolated_switch_large_0[3|2]/on avdd isolated_switch_large_0[3|2]/off
+ dvdd left_instramp_out ulpcomp_p dvss isolated_switch_large
Xisolated_switch_large_0[4|2] avss isolated_switch_large_0[4|2]/on avdd isolated_switch_large_0[4|2]/off
+ dvdd left_instramp_out comp_p dvss isolated_switch_large
Xisolated_switch_large_0[5|2] avss isolated_switch_large_0[5|2]/on avdd isolated_switch_large_0[5|2]/off
+ dvdd left_instramp_out adc0 dvss isolated_switch_large
.ends

.subckt audiodac_drv_latch in_p in_n vdd_hi vss
X0 in_p in_n vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X1 vss in_p in_n vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X2 in_n in_p vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X3 vdd_hi in_n in_p vdd_hi sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X4 in_p in_n vdd_hi vdd_hi sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X5 vdd_hi in_p in_n vdd_hi sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X6 in_n in_p vdd_hi vdd_hi sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X7 vss in_n in_p vss sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CYU746 a_n503_n1000# a_n345_n1000# a_n819_n1000#
+ a_29_n1097# a_n187_n1000# a_n661_n1000# a_n129_n1097# a_n603_n1097# w_n1019_n1297#
+ a_503_n1097# a_n445_n1097# a_345_n1097# a_n287_n1097# a_187_n1097# a_n761_n1097#
+ a_129_n1000# a_661_n1097# a_603_n1000# a_445_n1000# a_287_n1000# a_761_n1000# a_n29_n1000#
X0 a_445_n1000# a_345_n1097# a_287_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X1 a_n503_n1000# a_n603_n1097# a_n661_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X2 a_n29_n1000# a_n129_n1097# a_n187_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X3 a_603_n1000# a_503_n1097# a_445_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X4 a_n661_n1000# a_n761_n1097# a_n819_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X5 a_n187_n1000# a_n287_n1097# a_n345_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X6 a_761_n1000# a_661_n1097# a_603_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X7 a_287_n1000# a_187_n1097# a_129_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X8 a_n345_n1000# a_n445_n1097# a_n503_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X9 a_129_n1000# a_29_n1097# a_n29_n1000# w_n1019_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_QABAEG a_30_n588# a_288_n500# a_n478_n722# a_n128_n588#
+ a_188_n588# a_n286_n588# a_130_n500# a_n28_n500# a_n186_n500# a_n344_n500#
X0 a_n28_n500# a_n128_n588# a_n186_n500# a_n478_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X1 a_288_n500# a_188_n588# a_130_n500# a_n478_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X2 a_n186_n500# a_n286_n588# a_n344_n500# a_n478_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X3 a_130_n500# a_30_n588# a_n28_n500# a_n478_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3__0 a_n242_n622# a_50_n400# a_n108_n400#
+ a_n50_n488#
X0 a_50_n400# a_n50_n488# a_n108_n400# a_n242_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_YSH3F7 a_503_n1088# a_n445_n1088# a_n953_n1222#
+ a_n503_n1000# a_345_n1088# a_n287_n1088# a_n345_n1000# a_n819_n1000# a_187_n1088#
+ a_n761_n1088# a_n187_n1000# a_661_n1088# a_n661_n1000# a_129_n1000# a_29_n1088#
+ a_603_n1000# a_445_n1000# a_287_n1000# a_n129_n1088# a_761_n1000# a_n29_n1000# a_n603_n1088#
X0 a_n503_n1000# a_n603_n1088# a_n661_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X1 a_n29_n1000# a_n129_n1088# a_n187_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X2 a_603_n1000# a_503_n1088# a_445_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X3 a_n661_n1000# a_n761_n1088# a_n819_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X4 a_n187_n1000# a_n287_n1088# a_n345_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X5 a_761_n1000# a_661_n1088# a_603_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X6 a_287_n1000# a_187_n1088# a_129_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X7 a_n345_n1000# a_n445_n1088# a_n503_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X8 a_129_n1000# a_29_n1088# a_n29_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X9 a_445_n1000# a_345_n1088# a_287_n1000# a_n953_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_QCNVDG a_n108_n1000# a_n366_n1088# a_n424_n1000#
+ a_266_n1088# a_n266_n1000# a_50_n1000# a_208_n1000# a_366_n1000# a_n50_n1088# a_n208_n1088#
+ a_108_n1088# a_n558_n1222#
X0 a_n266_n1000# a_n366_n1088# a_n424_n1000# a_n558_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X1 a_366_n1000# a_266_n1088# a_208_n1000# a_n558_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X2 a_50_n1000# a_n50_n1088# a_n108_n1000# a_n558_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X3 a_n108_n1000# a_n208_n1088# a_n266_n1000# a_n558_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X4 a_208_n1000# a_108_n1088# a_50_n1000# a_n558_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_WECJAU a_30_n1098# a_n28_n1000# a_n344_n1000#
+ a_n186_n1000# a_130_n1000# a_188_n1098# a_n128_n1098# a_288_n1000# a_n286_n1098#
+ w_n544_n1296#
X0 a_n28_n1000# a_n128_n1098# a_n186_n1000# w_n544_n1296# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X1 a_288_n1000# a_188_n1098# a_130_n1000# w_n544_n1296# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X2 a_n186_n1000# a_n286_n1098# a_n344_n1000# w_n544_n1296# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X3 a_130_n1000# a_30_n1098# a_n28_n1000# w_n544_n1296# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_54K6JW a_445_118# a_n345_118# a_n661_n2118# a_n187_118#
+ a_187_21# a_287_118# a_n445_21# a_n819_118# a_n661_118# a_761_118# a_345_21# a_29_21#
+ a_n603_21# a_129_n2118# a_29_n2215# a_603_n2118# a_503_21# a_445_n2118# a_287_n2118#
+ a_n129_n2215# a_761_n2118# a_n29_n2118# a_129_118# a_n129_21# a_n761_21# a_n603_n2215#
+ w_n1019_n2415# a_503_n2215# a_n445_n2215# a_n29_118# a_661_21# a_n503_n2118# a_345_n2215#
+ a_n287_n2215# a_603_118# a_n503_118# a_n345_n2118# a_187_n2215# a_n761_n2215# a_n819_n2118#
+ a_n187_n2118# a_661_n2215# a_n287_21#
X0 a_n661_n2118# a_n761_n2215# a_n819_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X1 a_n29_n2118# a_n129_n2215# a_n187_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X2 a_n187_n2118# a_n287_n2215# a_n345_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X3 a_129_n2118# a_29_n2215# a_n29_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X4 a_n661_118# a_n761_21# a_n819_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X5 a_445_n2118# a_345_n2215# a_287_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X6 a_129_118# a_29_21# a_n29_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X7 a_n187_118# a_n287_21# a_n345_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X8 a_n345_118# a_n445_21# a_n503_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X9 a_n503_118# a_n603_21# a_n661_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X10 a_n345_n2118# a_n445_n2215# a_n503_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X11 a_n29_118# a_n129_21# a_n187_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X12 a_603_n2118# a_503_n2215# a_445_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X13 a_761_118# a_661_21# a_603_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X14 a_761_n2118# a_661_n2215# a_603_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X15 a_287_118# a_187_21# a_129_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X16 a_445_118# a_345_21# a_287_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X17 a_n503_n2118# a_n603_n2215# a_n661_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X18 a_603_118# a_503_21# a_445_118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X19 a_287_n2118# a_187_n2215# a_129_n2118# w_n1019_n2415# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_HKUKAU a_30_n162# w_n386_n362# a_n28_n64# a_n128_n162#
+ a_n186_n64# a_130_n64#
X0 a_n28_n64# a_n128_n162# a_n186_n64# w_n386_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X1 a_130_n64# a_30_n162# a_n28_n64# w_n386_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3QQKN5 a_130_n400# w_n386_n696# a_n28_n400# a_n186_n400#
+ a_n128_n498# a_30_n498#
X0 a_n28_n400# a_n128_n498# a_n186_n400# w_n386_n696# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_130_n400# a_30_n498# a_n28_n400# w_n386_n696# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt audiodac_drv_lite_half in crosscon out vdd_hi vss
Xsky130_fd_pr__pfet_g5v0d10v5_CYU746_0 vdd_hi drv4 vdd_hi crosscon vdd_hi drv4 crosscon
+ crosscon vdd_hi crosscon crosscon crosscon crosscon crosscon crosscon vdd_hi crosscon
+ drv4 vdd_hi drv4 vdd_hi drv4 sky130_fd_pr__pfet_g5v0d10v5_CYU746
Xsky130_fd_pr__nfet_g5v0d10v5_QABAEG_0 drv2 vss vss drv2 drv2 drv2 crosscon vss crosscon
+ vss sky130_fd_pr__nfet_g5v0d10v5_QABAEG
Xsky130_fd_pr__nfet_g5v0d10v5_MJGQJ3_0 vss drv2 vss drv1 sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3__0
Xsky130_fd_pr__nfet_g5v0d10v5_RX3AJQ_0 vss vss drv1 in sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ
Xsky130_fd_pr__nfet_g5v0d10v5_YSH3F7_0 drv4 drv4 vss vss drv4 drv4 out vss drv4 drv4
+ vss drv4 out vss drv4 out vss out drv4 vss out drv4 sky130_fd_pr__nfet_g5v0d10v5_YSH3F7
Xsky130_fd_pr__nfet_g5v0d10v5_YSH3F7_1 drv4 drv4 vss vss drv4 drv4 out vss drv4 drv4
+ vss drv4 out vss drv4 out vss out drv4 vss out drv4 sky130_fd_pr__nfet_g5v0d10v5_YSH3F7
Xsky130_fd_pr__nfet_g5v0d10v5_QCNVDG_0 vss crosscon vss crosscon drv4 drv4 vss drv4
+ crosscon crosscon crosscon vss sky130_fd_pr__nfet_g5v0d10v5_QCNVDG
Xsky130_fd_pr__pfet_g5v0d10v5_WECJAU_0 drv2 vdd_hi vdd_hi crosscon crosscon drv2 drv2
+ vdd_hi drv2 vdd_hi sky130_fd_pr__pfet_g5v0d10v5_WECJAU
Xsky130_fd_pr__pfet_g5v0d10v5_54K6JW_0 vdd_hi out out vdd_hi drv4 out drv4 vdd_hi
+ out vdd_hi drv4 drv4 drv4 vdd_hi drv4 out drv4 vdd_hi out drv4 vdd_hi out vdd_hi
+ drv4 drv4 drv4 vdd_hi drv4 drv4 out drv4 vdd_hi drv4 drv4 out vdd_hi out drv4 drv4
+ vdd_hi vdd_hi drv4 drv4 sky130_fd_pr__pfet_g5v0d10v5_54K6JW
Xsky130_fd_pr__pfet_g5v0d10v5_54K6JW_1 vdd_hi out out vdd_hi drv4 out drv4 vdd_hi
+ out vdd_hi drv4 drv4 drv4 vdd_hi drv4 out drv4 vdd_hi out drv4 vdd_hi out vdd_hi
+ drv4 drv4 drv4 vdd_hi drv4 drv4 out drv4 vdd_hi drv4 drv4 out vdd_hi out drv4 drv4
+ vdd_hi vdd_hi drv4 drv4 sky130_fd_pr__pfet_g5v0d10v5_54K6JW
Xsky130_fd_pr__pfet_g5v0d10v5_HKUKAU_0 in vdd_hi vdd_hi in drv1 drv1 sky130_fd_pr__pfet_g5v0d10v5_HKUKAU
Xsky130_fd_pr__pfet_g5v0d10v5_3QQKN5_1 vdd_hi vdd_hi drv2 vdd_hi drv1 drv1 sky130_fd_pr__pfet_g5v0d10v5_3QQKN5
.ends

.subckt sky130_fd_pr__nfet_01v8_U85QGS a_62_n200# a_n368_222# a_n224_n200# a_n320_n200#
+ a_398_222# a_n32_n200# a_n508_n200# a_302_n288# a_14_222# a_n464_n288# a_446_n200#
+ a_206_222# a_158_n200# a_110_n288# a_n272_n288# a_254_n200# a_n610_n374# a_n176_222#
+ a_350_n200# a_n416_n200# a_n128_n200# a_n80_n288#
X0 a_n128_n200# a_n176_222# a_n224_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1 a_n416_n200# a_n464_n288# a_n508_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2 a_n320_n200# a_n368_222# a_n416_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3 a_n32_n200# a_n80_n288# a_n128_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.32 pd=2.32 as=0.33 ps=2.33 w=2 l=0.15
X4 a_350_n200# a_302_n288# a_254_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X5 a_254_n200# a_206_222# a_158_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X6 a_158_n200# a_110_n288# a_62_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X7 a_n224_n200# a_n272_n288# a_n320_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X8 a_446_n200# a_398_222# a_350_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X9 a_62_n200# a_14_222# a_n32_n200# a_n610_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.32 ps=2.32 w=2 l=0.15
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_B24TY6 a_n50_n298# a_50_n200# a_n108_n200# a_n266_n200#
+ w_n624_n496# a_n424_n200# a_108_n298# a_n208_n298# a_266_n298# a_208_n200# a_n366_n298#
+ a_366_n200#
X0 a_n108_n200# a_n208_n298# a_n266_n200# w_n624_n496# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X1 a_208_n200# a_108_n298# a_50_n200# w_n624_n496# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X2 a_n266_n200# a_n366_n298# a_n424_n200# w_n624_n496# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X3 a_366_n200# a_266_n298# a_208_n200# w_n624_n496# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X4 a_50_n200# a_n50_n298# a_n108_n200# w_n624_n496# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_ARHMTT a_n148_n1000# a_n386_n1000# a_566_n1000#
+ a_328_n1000# a_90_n1000# a_n758_n1222# a_n566_n1088# a_n328_n1088# a_n624_n1000#
+ a_n90_n1088# a_386_n1088# a_148_n1088#
X0 a_n148_n1000# a_n328_n1088# a_n386_n1000# a_n758_n1222# sky130_fd_pr__nfet_05v0_nvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.9
X1 a_90_n1000# a_n90_n1088# a_n148_n1000# a_n758_n1222# sky130_fd_pr__nfet_05v0_nvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.9
X2 a_566_n1000# a_386_n1088# a_328_n1000# a_n758_n1222# sky130_fd_pr__nfet_05v0_nvt ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.9
X3 a_328_n1000# a_148_n1088# a_90_n1000# a_n758_n1222# sky130_fd_pr__nfet_05v0_nvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.9
X4 a_n386_n1000# a_n566_n1088# a_n624_n1000# a_n758_n1222# sky130_fd_pr__nfet_05v0_nvt ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.9
.ends

.subckt audiodac_drv_ls in_p in_n out_p out_n vdd_hi vdd_lo VSUBS
XXM1 VSUBS in_p a_n3307_n18881# VSUBS in_p a_n3307_n18881# VSUBS in_p in_p in_p VSUBS
+ in_p a_n3307_n18881# in_p in_p VSUBS VSUBS in_p a_n3307_n18881# a_n3307_n18881#
+ VSUBS in_p sky130_fd_pr__nfet_01v8_U85QGS
XXM5 out_n vdd_hi out_p vdd_hi vdd_hi out_p out_n out_n out_n out_p out_n vdd_hi sky130_fd_pr__pfet_g5v0d10v5_B24TY6
XXM6 out_p vdd_hi out_n vdd_hi vdd_hi out_n out_p out_p out_p out_n out_p vdd_hi sky130_fd_pr__pfet_g5v0d10v5_B24TY6
Xsky130_fd_pr__nfet_05v0_nvt_ARHMTT_0 out_n a_n3307_n18881# a_n3307_n18881# out_n
+ a_n3307_n18881# VSUBS vdd_lo vdd_lo out_n vdd_lo vdd_lo vdd_lo sky130_fd_pr__nfet_05v0_nvt_ARHMTT
Xsky130_fd_pr__nfet_01v8_U85QGS_0 VSUBS in_n m1_n1994_n18882# VSUBS in_n m1_n1994_n18882#
+ VSUBS in_n in_n in_n VSUBS in_n m1_n1994_n18882# in_n in_n VSUBS VSUBS in_n m1_n1994_n18882#
+ m1_n1994_n18882# VSUBS in_n sky130_fd_pr__nfet_01v8_U85QGS
Xsky130_fd_pr__nfet_05v0_nvt_ARHMTT_1 m1_n1994_n18882# out_p out_p m1_n1994_n18882#
+ out_p VSUBS vdd_lo vdd_lo m1_n1994_n18882# vdd_lo vdd_lo vdd_lo sky130_fd_pr__nfet_05v0_nvt_ARHMTT
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_VDASXE a_n1058_n5500# a_n1000_n5597# w_n1258_n5797#
+ a_1000_n5500#
X0 a_1000_n5500# a_n1000_n5597# a_n1058_n5500# w_n1258_n5797# sky130_fd_pr__pfet_g5v0d10v5 ad=15.95 pd=110.58 as=15.95 ps=110.58 w=55 l=10
.ends

.subckt sky130_iic_ip__audiodac_drv_lite in_p in_n out_p out_n in_hi vdd vss
Xaudiodac_drv_latch_0 audiodac_drv_latch_0/in_p audiodac_drv_latch_0/in_n vdd vss
+ audiodac_drv_latch
Xaudiodac_drv_lite_half_0 audiodac_drv_ls_0/out_n audiodac_drv_latch_0/in_n out_n
+ vdd vss audiodac_drv_lite_half
Xaudiodac_drv_lite_half_1 audiodac_drv_ls_0/out_p audiodac_drv_latch_0/in_p out_p
+ vdd vss audiodac_drv_lite_half
Xaudiodac_drv_ls_0 in_p in_n audiodac_drv_ls_0/out_p audiodac_drv_ls_0/out_n vdd in_hi
+ vss audiodac_drv_ls
Xsky130_fd_pr__pfet_g5v0d10v5_VDASXE_0 vdd vss vdd vdd sky130_fd_pr__pfet_g5v0d10v5_VDASXE
Xsky130_fd_pr__pfet_g5v0d10v5_VDASXE_1 vdd vss vdd vdd sky130_fd_pr__pfet_g5v0d10v5_VDASXE
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YHAZV5 a_n300_n197# a_300_n100# w_n558_n397#
+ a_n358_n100#
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n558_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_37RBXE a_n147_n172# a_n45_n70#
X0 a_n147_n172# a_n45_n70# sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EEVBR7 a_n300_n288# a_300_n200# a_n492_n422#
+ a_n358_n200#
X0 a_300_n200# a_n300_n288# a_n358_n200# a_n492_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
.ends

.subckt sky130_fd_pr__nfet_01v8_MG6U6H a_300_n100# a_n358_n100# a_n300_n188# a_n460_n274#
X0 a_300_n100# a_n300_n188# a_n358_n100# a_n460_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__pfet_01v8_J2L9Q3 a_n300_n197# a_300_n100# a_n358_n100# w_n496_n319#
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n496_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt ov_level_shifter in out out_b dvss avss dvdd avdd
Xsky130_fd_pr__pfet_g5v0d10v5_YHAZV5_0 out_b out avdd avdd sky130_fd_pr__pfet_g5v0d10v5_YHAZV5
Xsky130_fd_pr__pfet_g5v0d10v5_YHAZV5_1 out out_b avdd avdd sky130_fd_pr__pfet_g5v0d10v5_YHAZV5
Xsky130_fd_pr__diode_pw2nd_05v5_37RBXE_0 dvss in sky130_fd_pr__diode_pw2nd_05v5_37RBXE
Xsky130_fd_pr__nfet_g5v0d10v5_EEVBR7_0 in_b out avss avss sky130_fd_pr__nfet_g5v0d10v5_EEVBR7
Xsky130_fd_pr__nfet_g5v0d10v5_EEVBR7_1 in out_b avss avss sky130_fd_pr__nfet_g5v0d10v5_EEVBR7
Xsky130_fd_pr__nfet_01v8_MG6U6H_0 dvss in_b in dvss sky130_fd_pr__nfet_01v8_MG6U6H
Xsky130_fd_pr__pfet_01v8_J2L9Q3_0 in in_b dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9Q3
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_F6RBXN a_n147_n172# a_n45_n70#
X0 a_n147_n172# a_n45_n70# sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_6H9SQ3 a_n300_n197# a_300_n100# w_n558_n397#
+ a_n358_n100#
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n558_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CY564Z a_300_n100# a_n492_n322# a_n358_n100#
+ a_n300_n188#
X0 a_300_n100# a_n300_n188# a_n358_n100# a_n492_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt trans_gate_m in ena_b ena out avdd vss
Xsky130_fd_pr__pfet_g5v0d10v5_6H9SQ3_1 ena_b out avdd in sky130_fd_pr__pfet_g5v0d10v5_6H9SQ3
Xsky130_fd_pr__nfet_g5v0d10v5_CY564Z_0 out vss in ena sky130_fd_pr__nfet_g5v0d10v5_CY564Z
.ends

.subckt ov_multiplexer in_0000 in_0001 in_0010 in_0011 in_0100 in_0101 in_0110 in_0111
+ vtrip_3 vtrip_3_b vtrip_2 vtrip_1 out vtrip_1_b vtrip_0 vtrip_0_b in_1000 in_1001
+ in_1010 in_1011 in_1100 in_1101 in_1110 in_1111 vtrip_2_b avdd_uq0 avdd_uq3 avdd_uq1
+ avdd_uq2 vss avdd
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_2 vss vtrip_0_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_3 vss vtrip_0 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_4 vss vtrip_1 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_5 vss vtrip_1_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_6 vss vtrip_1_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_7 vss vtrip_1 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_8 vss vtrip_2_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_9 vss vtrip_2 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xtrans_gate_m_20 trans_gate_m_20/in vtrip_2 vtrip_2_b trans_gate_m_33/in avdd vss
+ trans_gate_m
Xtrans_gate_m_31 trans_gate_m_31/in vtrip_1 vtrip_1_b trans_gate_m_20/in avdd_uq1
+ vss trans_gate_m
Xtrans_gate_m_0 in_0010 vtrip_0 vtrip_0_b trans_gate_m_29/in avdd_uq2 vss trans_gate_m
Xtrans_gate_m_1 in_0011 vtrip_0_b vtrip_0 trans_gate_m_29/in avdd_uq2 vss trans_gate_m
Xtrans_gate_m_10 in_1000 vtrip_0 vtrip_0_b trans_gate_m_23/in avdd_uq3 vss trans_gate_m
Xtrans_gate_m_21 trans_gate_m_5/out vtrip_1_b vtrip_1 trans_gate_m_32/in avdd_uq1
+ vss trans_gate_m
Xtrans_gate_m_32 trans_gate_m_32/in vtrip_2 vtrip_2_b trans_gate_m_34/in avdd vss
+ trans_gate_m
Xtrans_gate_m_2 in_0110 vtrip_0 vtrip_0_b trans_gate_m_3/out avdd_uq2 vss trans_gate_m
Xtrans_gate_m_11 in_1001 vtrip_0_b vtrip_0 trans_gate_m_23/in avdd_uq3 vss trans_gate_m
Xtrans_gate_m_33 trans_gate_m_33/in vtrip_3 vtrip_3_b out avdd_uq0 vss trans_gate_m
Xtrans_gate_m_3 in_0111 vtrip_0_b vtrip_0 trans_gate_m_3/out avdd_uq2 vss trans_gate_m
Xtrans_gate_m_12 in_0101 vtrip_0_b vtrip_0 trans_gate_m_27/in avdd_uq3 vss trans_gate_m
Xtrans_gate_m_23 trans_gate_m_23/in vtrip_1 vtrip_1_b trans_gate_m_32/in avdd_uq1
+ vss trans_gate_m
Xtrans_gate_m_34 trans_gate_m_34/in vtrip_3_b vtrip_3 out avdd_uq0 vss trans_gate_m
Xtrans_gate_m_4 in_1011 vtrip_0_b vtrip_0 trans_gate_m_5/out avdd_uq2 vss trans_gate_m
Xtrans_gate_m_13 in_0100 vtrip_0 vtrip_0_b trans_gate_m_27/in avdd_uq3 vss trans_gate_m
Xtrans_gate_m_5 in_1010 vtrip_0 vtrip_0_b trans_gate_m_5/out avdd_uq2 vss trans_gate_m
Xtrans_gate_m_14 in_0001 vtrip_0_b vtrip_0 trans_gate_m_31/in avdd_uq3 vss trans_gate_m
Xtrans_gate_m_25 trans_gate_m_3/out vtrip_1_b vtrip_1 trans_gate_m_28/in avdd_uq1
+ vss trans_gate_m
Xtrans_gate_m_6 in_1110 vtrip_0 vtrip_0_b trans_gate_m_7/out avdd_uq2 vss trans_gate_m
Xtrans_gate_m_15 in_0000 vtrip_0 vtrip_0_b trans_gate_m_31/in avdd_uq3 vss trans_gate_m
Xtrans_gate_m_27 trans_gate_m_27/in vtrip_1 vtrip_1_b trans_gate_m_28/in avdd_uq1
+ vss trans_gate_m
Xtrans_gate_m_37 trans_gate_m_37/in vtrip_2_b vtrip_2 trans_gate_m_34/in avdd vss
+ trans_gate_m
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_10 vss vtrip_3_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xtrans_gate_m_7 in_1111 vtrip_0_b vtrip_0 trans_gate_m_7/out avdd_uq2 vss trans_gate_m
Xtrans_gate_m_28 trans_gate_m_28/in vtrip_2_b vtrip_2 trans_gate_m_33/in avdd vss
+ trans_gate_m
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_11 vss vtrip_3 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xtrans_gate_m_8 in_1101 vtrip_0_b vtrip_0 trans_gate_m_9/out avdd_uq3 vss trans_gate_m
Xtrans_gate_m_18 trans_gate_m_9/out vtrip_1 vtrip_1_b trans_gate_m_37/in avdd_uq1
+ vss trans_gate_m
Xtrans_gate_m_29 trans_gate_m_29/in vtrip_1_b vtrip_1 trans_gate_m_20/in avdd_uq1
+ vss trans_gate_m
Xtrans_gate_m_9 in_1100 vtrip_0 vtrip_0_b trans_gate_m_9/out avdd_uq3 vss trans_gate_m
Xtrans_gate_m_19 trans_gate_m_7/out vtrip_1_b vtrip_1 trans_gate_m_37/in avdd_uq1
+ vss trans_gate_m
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0 vss vtrip_0 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_1 vss vtrip_0_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_LV9PDH a_8742_125# a_n3732_n557# a_1560_125#
+ a_3828_n557# a_n7512_n557# a_804_n557# a_7608_n557# a_n4110_n557# a_3072_125# a_4206_n557#
+ a_4584_125# a_n4110_125# a_6096_125# a_n5622_125# a_6852_n557# a_n4866_n557# a_n1464_n557#
+ a_3450_n557# a_48_125# a_n8646_n557# a_7230_n557# a_n5244_n557# a_n7134_125# a_n8646_125#
+ a_n1464_125# a_n9024_n557# a_n2976_125# a_804_125# a_2316_125# a_3828_125# a_n7890_n557#
+ a_5340_125# a_7986_n557# a_n4488_125# a_4584_n557# a_n2598_n557# a_1182_n557# a_6852_125#
+ a_8364_n557# a_n6378_n557# a_8364_125# a_1182_125# a_2694_125# a_n2220_125# a_n1842_n557#
+ a_48_n557# a_1938_n557# a_n3732_125# a_n708_125# a_n5622_n557# a_n2220_n557# a_5718_n557#
+ a_2316_n557# a_6096_n557# a_n5244_125# a_n6000_n557# a_n6756_125# a_7608_125# a_n8268_125#
+ a_n2976_n557# a_4962_n557# a_n1086_125# a_1560_n557# a_1938_125# a_n2598_125# a_3450_125#
+ a_4962_125# a_8742_n557# a_5340_n557# a_n6756_n557# a_426_125# a_n3354_n557# a_6474_125#
+ a_n7134_n557# a_426_n557# a_7986_125# a_n708_n557# a_n6000_125# a_n7512_125# a_2694_n557#
+ a_n1842_125# a_6474_n557# a_3072_n557# a_n4488_n557# a_n1086_n557# a_n330_125# a_n9024_125#
+ a_n3354_125# a_n8268_n557# a_n4866_125# a_n330_n557# a_n7890_125# a_4206_125# a_5718_125#
+ a_7230_125# VSUBS a_n6378_125#
X0 a_n8646_125# a_n8646_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X1 a_n6000_125# a_n6000_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X2 a_n1464_125# a_n1464_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X3 a_6474_125# a_6474_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X4 a_804_125# a_804_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X5 a_n7134_125# a_n7134_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X6 a_n4488_125# a_n4488_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X7 a_5718_125# a_5718_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X8 a_6852_125# a_6852_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X9 a_n1842_125# a_n1842_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X10 a_n7512_125# a_n7512_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X11 a_n4866_125# a_n4866_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X12 a_4206_125# a_4206_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X13 a_5340_125# a_5340_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X14 a_n330_125# a_n330_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X15 a_2694_125# a_2694_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X16 a_n7890_125# a_n7890_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X17 a_n2220_125# a_n2220_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X18 a_n3354_125# a_n3354_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X19 a_8364_125# a_8364_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X20 a_n708_125# a_n708_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X21 a_1182_125# a_1182_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X22 a_1938_125# a_1938_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X23 a_n9024_125# a_n9024_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X24 a_48_125# a_48_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X25 a_n6378_125# a_n6378_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X26 a_n3732_125# a_n3732_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X27 a_7608_125# a_7608_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X28 a_8742_125# a_8742_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X29 a_1560_125# a_1560_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X30 a_n6756_125# a_n6756_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X31 a_7230_125# a_7230_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X32 a_4584_125# a_4584_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X33 a_n5244_125# a_n5244_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X34 a_n4110_125# a_n4110_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X35 a_n2598_125# a_n2598_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X36 a_3072_125# a_3072_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X37 a_3828_125# a_3828_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X38 a_4962_125# a_4962_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X39 a_n8268_125# a_n8268_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X40 a_n5622_125# a_n5622_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X41 a_n2976_125# a_n2976_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X42 a_n1086_125# a_n1086_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X43 a_6096_125# a_6096_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X44 a_7986_125# a_7986_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X45 a_426_125# a_426_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X46 a_2316_125# a_2316_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X47 a_3450_125# a_3450_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_H3F4MM a_1182_1930# a_n4488_n1826# a_7986_n1826#
+ a_n6378_n2362# a_n7890_5150# a_n7890_n5582# a_7986_5150# a_4584_5150# a_n2598_5150#
+ a_1182_5150# a_8364_1930# a_n6378_1930# a_n4866_n1826# a_n6756_n2362# a_8364_5150#
+ a_n6378_5150# a_n2598_n1826# a_n6000_n5582# a_n4488_n2362# a_n3732_1394# a_7986_n2362#
+ a_3828_1394# a_426_n5582# a_7230_n5582# a_7608_n5582# a_n2976_n1826# a_n4866_n2362#
+ a_n7512_1394# a_n4110_1394# a_804_1394# a_7608_1394# a_4206_1394# a_4206_n1826#
+ a_n1842_1930# a_n4110_n5582# a_804_n5582# a_n2598_n2362# a_48_1930# a_1938_1930#
+ a_5340_n5582# a_n1842_5150# a_5718_n5582# a_48_5150# a_1938_5150# a_n5622_1930#
+ a_n2976_n2362# a_n2220_1930# a_5718_1930# a_3072_n5582# a_2316_1930# a_n9024_n1826#
+ a_6096_1930# a_2316_n1826# a_4206_n2362# a_n2220_n5582# a_n5622_5150# a_n2220_5150#
+ a_5718_5150# a_2316_5150# a_6852_1394# a_n6000_1930# a_6096_5150# a_n4866_1394#
+ a_3450_1394# a_3450_n5582# a_3828_n5582# a_n1464_1394# a_n8268_n5582# a_n6000_5150#
+ a_1182_n5582# a_n7134_n1826# a_n9024_n2362# a_2316_n2362# a_n8646_1394# a_7230_1394#
+ a_n5244_1394# a_8364_n1826# a_4962_1930# a_n2976_1930# a_1560_1930# a_n8646_n5582#
+ a_1560_n5582# a_n7512_n1826# a_1938_n5582# a_6096_n1826# a_n9024_1394# a_4962_5150#
+ a_n2976_5150# a_n6378_n5582# a_n5244_n1826# a_n7134_n2362# a_1560_5150# a_8742_n1826#
+ a_8742_1930# a_n6756_1930# a_5340_1930# a_n3354_1930# a_n330_n1826# a_6474_n1826#
+ a_n708_n1826# a_8364_n2362# a_8742_5150# a_n6756_n5582# a_n6756_5150# a_n5622_n1826#
+ a_5340_5150# a_n7512_n2362# a_48_n1826# a_n7890_1394# a_n3354_5150# a_6096_n2362#
+ a_n7134_1930# a_7986_1394# a_n4488_n5582# a_426_1930# a_4584_1394# a_7986_n5582#
+ a_n3354_n1826# a_n2598_1394# a_6852_n1826# a_n5244_n2362# a_8742_n2362# a_1182_1394#
+ a_n708_1930# a_n7134_5150# a_n1086_n1826# a_426_5150# a_4584_n1826# a_n330_n2362#
+ a_6474_n2362# a_n708_n2362# a_8364_1394# a_n4866_n5582# a_n3732_n1826# a_n6378_1394#
+ a_n5622_n2362# a_48_n2362# a_n708_5150# a_2694_1930# a_n2598_n5582# a_n1464_n1826#
+ a_4962_n1826# a_n3354_n2362# a_6852_n2362# a_2694_5150# a_2694_n1826# a_n1086_n2362#
+ a_4584_n2362# a_6474_1930# a_n2976_n5582# a_n4488_1930# a_n1842_n1826# a_n3732_n2362#
+ a_3072_1930# a_n1086_1930# a_4206_n5582# a_6474_5150# a_n1464_n2362# a_4962_n2362#
+ a_n4488_5150# a_3072_5150# a_n1842_1394# a_n1086_5150# a_n8268_1930# a_48_1394#
+ a_1938_1394# a_2694_n2362# a_n330_1930# a_n1842_n2362# a_n8268_5150# a_n5622_1394#
+ a_n9024_n5582# a_n2220_1394# a_2316_n5582# a_5718_1394# a_n7890_n1826# a_n330_5150#
+ a_2316_1394# a_6096_1394# a_n6000_1394# a_n3732_1930# a_n7134_n5582# a_3828_1930#
+ a_n6000_n1826# a_n7890_n2362# a_n3732_5150# a_8364_n5582# a_426_n1826# a_7230_n1826#
+ a_3828_5150# a_7608_n1826# a_n7512_1930# a_n7512_n5582# a_n4110_1930# a_804_1930#
+ a_7608_1930# a_4962_1394# a_n2976_1394# a_4206_1930# a_1560_1394# a_6096_n5582#
+ a_n7512_5150# a_n5244_n5582# a_n4110_n1826# a_8742_n5582# a_804_n1826# a_n6000_n2362#
+ a_n4110_5150# a_804_5150# a_7608_5150# a_4206_5150# a_8742_1394# a_n6756_1394# a_5340_1394#
+ a_n3354_1394# a_6474_n5582# a_n330_n5582# a_n708_n5582# a_5340_n1826# a_426_n2362#
+ a_5718_n1826# a_7230_n2362# a_7608_n2362# a_n5622_n5582# a_48_n5582# a_3072_n1826#
+ a_n7134_1394# a_n3354_n5582# a_6852_n5582# a_n2220_n1826# a_n4110_n2362# a_804_n2362#
+ a_426_1394# a_6852_1930# a_n4866_1930# a_3450_1930# a_n1464_1930# a_n1086_n5582#
+ a_4584_n5582# a_n708_1394# a_3450_n1826# a_5340_n2362# a_3828_n1826# a_5718_n2362#
+ a_n3732_n5582# a_6852_5150# a_n4866_5150# a_3450_5150# a_n1464_5150# a_n8268_n1826#
+ a_1182_n1826# a_n8646_1930# a_3072_n2362# a_7230_1930# a_n5244_1930# a_n1464_n5582#
+ a_4962_n5582# a_n2220_n2362# a_2694_1394# a_n8646_5150# a_7230_5150# a_2694_n5582#
+ a_n8646_n1826# a_n5244_5150# a_1560_n1826# a_1938_n1826# a_3450_n2362# a_3828_n2362#
+ a_n9024_1930# a_n1842_n5582# a_6474_1394# a_n4488_1394# a_3072_1394# a_n6378_n1826#
+ a_n8268_n2362# a_n1086_1394# a_1182_n2362# a_n9024_5150# a_n8268_1394# a_n7890_1930#
+ a_n6756_n1826# a_n8646_n2362# a_1560_n2362# a_1938_n2362# a_7986_1930# VSUBS a_4584_1930#
+ a_n2598_1930# a_n330_1394#
X0 a_n1464_1394# a_n1464_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X1 a_n2598_n2362# a_n2598_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X2 a_4584_5150# a_4584_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X3 a_426_1394# a_426_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X4 a_n3732_1394# a_n3732_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X5 a_n4866_n2362# a_n4866_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X6 a_n1464_n2362# a_n1464_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X7 a_426_n2362# a_426_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X8 a_n3732_n2362# a_n3732_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X9 a_n5244_5150# a_n5244_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X10 a_n4110_5150# a_n4110_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X11 a_n2598_5150# a_n2598_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X12 a_3072_5150# a_3072_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X13 a_3828_5150# a_3828_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X14 a_4962_5150# a_4962_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X15 a_n9024_1394# a_n9024_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X16 a_6474_1394# a_6474_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X17 a_n8268_5150# a_n8268_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X18 a_n9024_n2362# a_n9024_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X19 a_8742_1394# a_8742_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X20 a_5718_1394# a_5718_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X21 a_n330_1394# a_n330_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X22 a_3072_1394# a_3072_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X23 a_n7890_1394# a_n7890_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X24 a_n5622_5150# a_n5622_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X25 a_n1086_5150# a_n1086_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X26 a_6096_5150# a_6096_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X27 a_6474_n2362# a_6474_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X28 a_5340_1394# a_5340_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X29 a_2316_1394# a_2316_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X30 a_8742_n2362# a_8742_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X31 a_5718_n2362# a_5718_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X32 a_n330_n2362# a_n330_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X33 a_n4488_1394# a_n4488_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X34 a_n2976_5150# a_n2976_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X35 a_7986_5150# a_7986_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X36 a_2316_5150# a_2316_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X37 a_3450_5150# a_3450_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X38 a_3072_n2362# a_3072_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X39 a_n6756_1394# a_n6756_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X40 a_426_5150# a_426_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X41 a_5340_n2362# a_5340_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X42 a_n7890_n2362# a_n7890_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X43 a_2316_n2362# a_2316_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X44 a_n1086_1394# a_n1086_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X45 a_n3354_1394# a_n3354_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X46 a_n4488_n2362# a_n4488_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X47 a_n5622_1394# a_n5622_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X48 a_n6756_n2362# a_n6756_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X49 a_n1086_n2362# a_n1086_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X50 a_n8646_5150# a_n8646_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X51 a_n3354_n2362# a_n3354_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X52 a_n5622_n2362# a_n5622_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X53 a_n6000_5150# a_n6000_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X54 a_n1464_5150# a_n1464_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X55 a_6474_5150# a_6474_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X56 a_804_5150# a_804_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X57 a_n7134_5150# a_n7134_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X58 a_6096_1394# a_6096_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X59 a_n4488_5150# a_n4488_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X60 a_8364_1394# a_8364_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X61 a_7608_1394# a_7608_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X62 a_5718_5150# a_5718_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X63 a_n1842_5150# a_n1842_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X64 a_6852_5150# a_6852_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X65 a_6096_n2362# a_6096_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X66 a_8364_n2362# a_8364_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X67 a_7230_1394# a_7230_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X68 a_4206_1394# a_4206_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X69 a_7608_n2362# a_7608_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X70 a_n6378_1394# a_n6378_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X71 a_n8646_1394# a_n8646_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X72 a_7230_n2362# a_7230_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X73 a_4206_n2362# a_4206_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X74 a_n5244_1394# a_n5244_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X75 a_n6378_n2362# a_n6378_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X76 a_n2220_1394# a_n2220_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X77 a_n7512_5150# a_n7512_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X78 a_n7512_1394# a_n7512_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X79 a_n8646_n2362# a_n8646_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X80 a_n4866_5150# a_n4866_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X81 a_2694_1394# a_2694_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X82 a_4206_5150# a_4206_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X83 a_n5244_n2362# a_n5244_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X84 a_4962_1394# a_4962_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X85 a_1938_1394# a_1938_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X86 a_5340_5150# a_5340_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X87 a_n2220_n2362# a_n2220_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X88 a_n7512_n2362# a_n7512_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X89 a_n330_5150# a_n330_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X90 a_2694_5150# a_2694_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X91 a_2694_n2362# a_2694_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X92 a_1560_1394# a_1560_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X93 a_48_1394# a_48_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X94 a_4962_n2362# a_4962_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X95 a_1938_n2362# a_1938_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X96 a_n2976_1394# a_n2976_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X97 a_1560_n2362# a_1560_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X98 a_48_n2362# a_48_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X99 a_n7890_5150# a_n7890_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X100 a_n1842_1394# a_n1842_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X101 a_n3354_5150# a_n3354_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X102 a_n2220_5150# a_n2220_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X103 a_8364_5150# a_8364_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X104 a_n2976_n2362# a_n2976_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X105 a_804_1394# a_804_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X106 a_1182_5150# a_1182_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X107 a_n1842_n2362# a_n1842_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X108 a_n708_5150# a_n708_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X109 a_1938_5150# a_1938_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X110 a_804_n2362# a_804_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X111 a_48_5150# a_48_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X112 a_n9024_5150# a_n9024_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X113 a_n8268_1394# a_n8268_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X114 a_n6378_5150# a_n6378_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X115 a_7608_5150# a_7608_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X116 a_n7134_1394# a_n7134_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X117 a_n3732_5150# a_n3732_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X118 a_8742_5150# a_8742_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X119 a_n8268_n2362# a_n8268_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X120 a_7986_1394# a_7986_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X121 a_n4110_1394# a_n4110_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X122 a_1560_5150# a_1560_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X123 a_4584_1394# a_4584_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X124 a_n7134_n2362# a_n7134_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X125 a_6852_1394# a_6852_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X126 a_3828_1394# a_3828_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X127 a_7986_n2362# a_7986_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X128 a_n4110_n2362# a_n4110_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X129 a_n708_1394# a_n708_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X130 a_1182_1394# a_1182_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X131 a_n6000_1394# a_n6000_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X132 a_4584_n2362# a_4584_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X133 a_3450_1394# a_3450_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X134 a_6852_n2362# a_6852_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X135 a_3828_n2362# a_3828_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X136 a_n2598_1394# a_n2598_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X137 a_n708_n2362# a_n708_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X138 a_n6756_5150# a_n6756_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X139 a_1182_n2362# a_1182_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X140 a_n4866_1394# a_n4866_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X141 a_3450_n2362# a_3450_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X142 a_n6000_n2362# a_n6000_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X143 a_7230_5150# a_7230_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_SB5CJ8 a_300_n300# a_n492_n522# a_n358_n300#
+ a_n300_n388#
X0 a_300_n300# a_n300_n388# a_n358_n300# a_n492_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=3
.ends

.subckt ov_voltage_divider avdd out_0000 out_0001 out_0010 out_0011 out_0100 out_0101
+ out_0110 out_0111 out_1000 out_1001 out_1010 out_1011 out_1100 out_1101 out_1110
+ out_1111 avss ena
Xsky130_fd_pr__res_xhigh_po_1p41_LV9PDH_0 avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss sky130_fd_pr__res_xhigh_po_1p41_LV9PDH
Xsky130_fd_pr__res_xhigh_po_1p41_LV9PDH_2 avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss sky130_fd_pr__res_xhigh_po_1p41_LV9PDH
Xsky130_fd_pr__res_xhigh_po_1p41_H3F4MM_0 m1_3399_9649# m1_7155_3979# m1_7155_16831#
+ m1_7155_2467# m1_179_955# m1_10911_577# m1_179_16831# m1_179_13051# m1_179_6247#
+ m1_179_10027# m1_3399_17209# m1_3399_2467# m1_7155_3979# m1_7155_2089# m1_179_16831#
+ m1_179_2467# m1_7155_6247# m1_10911_2845# out_1110 m1_3935_5113# m1_7155_16831#
+ m1_3935_12673# out_0011 m1_10911_15697# m1_10911_16453# m1_7155_5491# out_1110 m1_3399_1333#
+ m1_3935_4357# m1_3935_9649# m1_3935_16453# m1_3935_12673# m1_7155_13051# m1_3399_6625#
+ out_1101 out_0010 out_1000 m1_3399_8893# m1_3399_10405# m1_10911_14185# m1_179_7003#
+ m1_10911_14185# m1_179_8515# m1_179_10783# m1_3399_3223# out_1010 m1_3399_6625#
+ m1_3399_14185# m1_10911_11917# m1_3399_11161# avss m1_3399_14941# m1_7155_10783#
+ m1_7691_13051# out_0111 m1_179_3223# m1_179_6247# m1_179_14563# m1_179_10783# m1_3935_15697#
+ m1_3399_2845# m1_179_14563# m1_3399_3979# m1_3935_11917# m1_10911_11917# m1_10911_12673#
+ m1_3935_7381# m1_10911_577# m1_179_2467# out_0010 m1_7155_1711# avss m1_7691_10783#
+ m1_3399_199# m1_3935_15697# m1_3399_3601# m1_7155_17209# m1_3399_13429# m1_3399_5869#
+ m1_3399_10405# m1_10901_199# out_0001 m1_7155_1333# out_0001 m1_7155_14563# avss
+ m1_179_13807# m1_179_5491# m1_10911_2089# m1_7155_3601# m1_7155_1711# m1_179_10027#
+ avss avss m1_3399_2089# m1_3399_14185# m1_3399_5113# m1_7155_8515# m1_7155_15319#
+ m1_7155_7759# m1_7155_17209# avss m1_10911_2089# m1_179_1711# m1_7155_3223# m1_179_13807#
+ m1_7155_1333# m1_7155_8515# m1_3399_955# m1_179_5491# m1_7691_14563# m1_3399_1711#
+ m1_3935_16453# out_1101 m1_3399_8893# m1_3935_13429# m1_10911_16453# m1_7155_5491#
+ m1_3935_5869# m1_7155_15319# m1_7155_3601# avss m1_3935_9649# m1_3399_8137# m1_179_1711#
+ m1_7155_7759# m1_179_9271# m1_7155_13051# out_0100 m1_7691_15319# out_0101 m1_3399_17209#
+ out_1111 m1_7155_4735# m1_3399_2467# m1_7155_3223# out_0100 m1_179_7759# m1_3399_11161#
+ out_1001 m1_7155_7003# m1_7155_13807# out_1010 m1_7691_15319# m1_179_11539# m1_7155_11539#
+ out_0101 m1_7691_13051# m1_3399_14941# out_1001 m1_3399_4357# m1_7155_7003# out_1100
+ m1_3399_11917# m1_3399_7381# m1_10911_12673# m1_179_15319# m1_7691_7003# m1_7691_13807#
+ m1_179_3979# m1_179_11539# m1_3935_6625# m1_179_7759# m1_3399_577# m1_3935_8893#
+ m1_3935_10405# 51 m1_3399_8137# m1_7691_7003# m1_179_199# m1_3399_3223# avss m1_3935_6625#
+ out_0000 m1_3935_14185# m1_7155_955# m1_179_8515# m1_3935_11161# m1_3935_14941#
+ m1_3399_2845# m1_3399_5113# m1_10911_1333# m1_3399_12673# m1_7155_2845# m1_7155_955#
+ m1_179_4735# avdd m1_7155_9271# m1_7155_16075# m1_179_12295# m1_7155_16075# m1_3399_1333#
+ m1_10911_1333# m1_3399_4357# m1_3399_9649# m1_3399_16453# m1_3935_13429# m1_3935_5869#
+ m1_3399_12673# m1_3935_10405# m1_10911_14941# m1_179_955# out_1111 m1_7155_4735#
+ avss m1_7155_9271# m1_7155_2845# m1_179_4735# m1_179_9271# m1_179_16075# m1_179_13051#
+ avss m1_3399_2089# m1_3935_14185# m1_3935_5113# m1_10911_14941# m1_10901_8137# m1_10901_8137#
+ m1_7155_13807# m1_7691_9271# m1_7155_14563# m1_7691_16075# m1_7691_16075# m1_10911_2845#
+ out_0011 m1_7155_11539# m1_3399_1711# out_1011 m1_10911_15697# m1_7155_6247# out_1100
+ m1_7691_9271# m1_3935_8893# m1_3399_15697# m1_3399_3979# m1_3399_11917# m1_3399_7381#
+ out_0110 m1_10911_13429# m1_3935_8137# m1_7155_12295# m1_7691_13807# m1_7155_12295#
+ m1_7691_14563# out_1011 m1_179_15319# m1_179_3979# m1_179_12295# m1_179_7003# m1_7155_577#
+ m1_7155_10027# m1_3399_199# 51 m1_3399_15697# m1_3399_3601# out_0110 m1_10911_13429#
+ out_1000 m1_3935_11161# m1_179_199# m1_179_16075# out_0000 m1_7155_199# m1_179_3223#
+ m1_7155_10027# m1_7155_10783# m1_7691_12295# m1_7691_12295# avss out_0111 m1_3935_14941#
+ m1_3935_4357# m1_3935_11917# m1_7155_2467# m1_7155_577# m1_3935_7381# m1_7691_10027#
+ avss m1_3399_577# m1_3399_955# m1_7155_2089# m1_7155_199# m1_7691_10027# m1_7691_10783#
+ m1_3399_16453# avss m1_3399_13429# m1_3399_5869# m1_3935_8137# sky130_fd_pr__res_xhigh_po_1p41_H3F4MM
Xsky130_fd_pr__nfet_g5v0d10v5_SB5CJ8_0 avss avss m1_10901_199# ena sky130_fd_pr__nfet_g5v0d10v5_SB5CJ8
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0 avss ena sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
.ends

.subckt sky130_fd_pr__pfet_01v8_XTWSDC a_n1600_n197# a_1600_n100# a_n1658_n100# w_n1796_n319#
X0 a_1600_n100# a_n1600_n197# a_n1658_n100# w_n1796_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
.ends

.subckt sky130_fd_pr__nfet_01v8_7ZF23Z a_2000_n100# a_n2058_n100# a_n2000_n188# a_n2160_n274#
X0 a_2000_n100# a_n2000_n188# a_n2058_n100# a_n2160_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
.ends

.subckt sky130_fd_pr__nfet_01v8_V433WY a_300_n100# a_n358_n100# a_n300_n188# a_n460_n274#
X0 a_300_n100# a_n300_n188# a_n358_n100# a_n460_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_69BJMM a_n500_n188# a_500_n100# a_n692_n322#
+ a_n558_n100#
X0 a_500_n100# a_n500_n188# a_n558_n100# a_n692_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_E7V9VM w_n758_n897# a_n558_n600# a_n500_n697#
+ a_500_n600#
X0 a_500_n600# a_n500_n697# a_n558_n600# w_n758_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=5
.ends

.subckt trans_gate in ena_b ena out vss avdd
XXM1 ena out vss in sky130_fd_pr__nfet_g5v0d10v5_69BJMM
XXM2 avdd out ena_b in sky130_fd_pr__pfet_g5v0d10v5_E7V9VM
.ends

.subckt sky130_fd_pr__pfet_01v8_C2YSV5 a_n300_n197# a_300_n100# a_n358_n100# w_n496_n319#
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n496_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__pfet_01v8_J2L9E5 w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_GGMWVD w_n996_n319# a_n800_n197# a_800_n100# a_n858_n100#
X0 a_800_n100# a_n800_n197# a_n858_n100# w_n996_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
.ends

.subckt sky130_fd_pr__pfet_01v8_CDT3CS a_n1600_n197# a_1600_n100# a_n1658_n100# w_n1796_n319#
X0 a_1600_n100# a_n1600_n197# a_n1658_n100# w_n1796_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z a_100_n100# a_n292_n322# a_n158_n100#
+ a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n292_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_3HBZVM a_n158_n300# w_n296_n519# a_n100_n397# a_100_n300#
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n296_n519# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_697RXD a_800_n100# a_n858_n100# a_n800_n188# a_n960_n274#
X0 a_800_n100# a_n800_n188# a_n858_n100# a_n960_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_4T6WVE a_100_n130# a_n292_n352# a_n158_n130#
+ a_n100_n218#
X0 a_100_n130# a_n100_n218# a_n158_n130# a_n292_n352# sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_6975WM a_800_n130# a_n992_n352# a_n858_n130#
+ a_n800_n218#
X0 a_800_n130# a_n800_n218# a_n858_n130# a_n992_n352# sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DEN7YK a_800_n100# a_n992_n322# a_n858_n100#
+ a_n800_n188#
X0 a_800_n100# a_n800_n188# a_n858_n100# a_n992_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
.ends

.subckt sky130_fd_pr__pfet_01v8_G3L97A w_n996_n319# a_n800_n197# a_800_n100# a_n858_n100#
X0 a_800_n100# a_n800_n197# a_n858_n100# w_n996_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
.ends

.subckt sky130_fd_pr__nfet_01v8_C8TQ3N a_n158_n300# a_n100_n388# a_n260_n474# a_100_n300#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n260_n474# sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt comp_hyst out vref vin ena ibias dvss dvdd
XXMD16[0] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM12 dvss net1 net5 dvss sky130_fd_pr__nfet_01v8_7ZF23Z
XXM14 dvss net2 ena_b dvss sky130_fd_pr__nfet_01v8_V433WY
XXM13 dvss net5 ena_b dvss sky130_fd_pr__nfet_01v8_V433WY
Xx1 ibias ena_b ena net5 dvss dvdd trans_gate
XXM15 ena net4 dvdd dvdd sky130_fd_pr__pfet_01v8_C2YSV5
XXM16 ena net3 dvdd dvdd sky130_fd_pr__pfet_01v8_C2YSV5
XXM17 dvss out ena_b dvss sky130_fd_pr__nfet_01v8_V433WY
XXMD1[19] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM18 ena ena_b dvdd dvdd sky130_fd_pr__pfet_01v8_C2YSV5
XXMD1[18] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM19 dvss ena_b ena dvss sky130_fd_pr__nfet_01v8_V433WY
XXM6[3] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM3[1] dvdd net4 net4 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XXMD1[17] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM6[2] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8_CDT3CS
XXM3[0] dvdd net4 net4 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XXMD1[16] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM6[1] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM6[0] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8_CDT3CS
XXMD1[15] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[13] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[14] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[3] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[9] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[12] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[2] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[8] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[11] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[7] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[10] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[6] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[4] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[5] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XD1 dvss vref sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
XXMD1[3] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM7 dvdd net4 net2 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XD3 dvss ena sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
XXMD1[2] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM9 dvdd dvdd net3 out sky130_fd_pr__pfet_01v8_3HBZVM
XXM8 dvss net2 net2 dvss sky130_fd_pr__nfet_01v8_697RXD
XXMDN13[7] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXM1[1] net1 dvss net4 vref sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXMD1[1] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM1[0] net1 dvss net4 vref sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXM4[1] net3 net3 dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXMDN13[6] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMD1[0] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM4[0] net3 net3 dvdd dvdd sky130_fd_pr__pfet_01v8_CDT3CS
XXMDN13[5] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[4] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[3] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[2] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN8[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_DEN7YK
XXMDN8[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_DEN7YK
XXMD16[5] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXMD16[4] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM2[1] net1 dvss net3 vin sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXM5[1] dvdd net4 net3 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XXMD16[3] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM2[0] net1 dvss net3 vin sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXM5[0] dvdd net4 net3 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XXMD16[2] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXMD8[1] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_G3L97A
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0 dvss vin sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
XXM10 out net2 dvss dvss sky130_fd_pr__nfet_01v8_C8TQ3N
XXMD8[0] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_G3L97A
XXMD16[1] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM11 dvss net5 net5 dvss sky130_fd_pr__nfet_01v8_7ZF23Z
.ends

.subckt sky130_vbl_ip__overvoltage avdd dvdd ena vtrip[3] ibias vtrip[2] ovout vbg
+ vtrip[1] vtrip[0] dvss avss
Xov_level_shifter_0 vtrip[0] ov_level_shifter_0/out ov_level_shifter_0/out_b dvss
+ avss dvdd avdd ov_level_shifter
Xov_level_shifter_1 vtrip[1] ov_level_shifter_1/out ov_level_shifter_1/out_b dvss
+ avss dvdd avdd ov_level_shifter
Xov_level_shifter_2 vtrip[2] ov_level_shifter_2/out ov_level_shifter_2/out_b dvss
+ avss dvdd avdd ov_level_shifter
Xov_level_shifter_3 vtrip[3] ov_level_shifter_3/out ov_level_shifter_3/out_b dvss
+ avss dvdd avdd ov_level_shifter
Xov_multiplexer_0 ov_multiplexer_0/in_0000 ov_multiplexer_0/in_0001 ov_multiplexer_0/in_0010
+ ov_multiplexer_0/in_0011 ov_multiplexer_0/in_0100 ov_multiplexer_0/in_0101 ov_multiplexer_0/in_0110
+ ov_multiplexer_0/in_0111 ov_level_shifter_3/out ov_level_shifter_3/out_b ov_level_shifter_2/out
+ ov_level_shifter_1/out vin ov_level_shifter_1/out_b ov_level_shifter_0/out ov_level_shifter_0/out_b
+ ov_multiplexer_0/in_1000 ov_multiplexer_0/in_1001 ov_multiplexer_0/in_1010 ov_multiplexer_0/in_1011
+ ov_multiplexer_0/in_1100 ov_multiplexer_0/in_1101 ov_multiplexer_0/in_1110 ov_multiplexer_0/in_1111
+ ov_level_shifter_2/out_b avdd avdd avdd avdd avss avdd ov_multiplexer
Xov_voltage_divider_0 avdd ov_multiplexer_0/in_0000 ov_multiplexer_0/in_0001 ov_multiplexer_0/in_0010
+ ov_multiplexer_0/in_0011 ov_multiplexer_0/in_0100 ov_multiplexer_0/in_0101 ov_multiplexer_0/in_0110
+ ov_multiplexer_0/in_0111 ov_multiplexer_0/in_1000 ov_multiplexer_0/in_1001 ov_multiplexer_0/in_1010
+ ov_multiplexer_0/in_1011 ov_multiplexer_0/in_1100 ov_multiplexer_0/in_1101 ov_multiplexer_0/in_1110
+ ov_multiplexer_0/in_1111 avss ena ov_voltage_divider
Xcomp_hyst_0 ovout vbg vin ena ibias dvss dvdd comp_hyst
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_F5JQJ7 a_n445_n1088# a_n503_n1000# a_345_n1088#
+ a_n287_n1088# a_n345_n1000# a_187_n1088# a_n187_n1000# a_129_n1000# a_29_n1088#
+ a_445_n1000# a_287_n1000# a_n129_n1088# a_n637_n1222# a_n29_n1000#
X0 a_n29_n1000# a_n129_n1088# a_n187_n1000# a_n637_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X1 a_n187_n1000# a_n287_n1088# a_n345_n1000# a_n637_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X2 a_287_n1000# a_187_n1088# a_129_n1000# a_n637_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X3 a_n345_n1000# a_n445_n1088# a_n503_n1000# a_n637_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X4 a_129_n1000# a_29_n1088# a_n29_n1000# a_n637_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X5 a_445_n1000# a_345_n1088# a_287_n1000# a_n637_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AQSWZU a_n503_n1000# a_n345_n1000# a_n819_n1000#
+ a_29_n1097# a_n187_n1000# a_n661_n1000# a_n977_n1000# a_n129_n1097# a_n603_n1097#
+ a_503_n1097# a_n445_n1097# a_n919_n1097# a_345_n1097# a_n287_n1097# a_819_n1097#
+ a_187_n1097# a_n761_n1097# w_n1177_n1297# a_129_n1000# a_661_n1097# a_603_n1000#
+ a_919_n1000# a_445_n1000# a_287_n1000# a_761_n1000# a_n29_n1000#
X0 a_445_n1000# a_345_n1097# a_287_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X1 a_n503_n1000# a_n603_n1097# a_n661_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X2 a_n29_n1000# a_n129_n1097# a_n187_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X3 a_603_n1000# a_503_n1097# a_445_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X4 a_n819_n1000# a_n919_n1097# a_n977_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.5
X5 a_n661_n1000# a_n761_n1097# a_n819_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X6 a_919_n1000# a_819_n1097# a_761_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.5
X7 a_n187_n1000# a_n287_n1097# a_n345_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X8 a_761_n1000# a_661_n1097# a_603_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X9 a_287_n1000# a_187_n1097# a_129_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X10 a_n345_n1000# a_n445_n1097# a_n503_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
X11 a_129_n1000# a_29_n1097# a_n29_n1000# w_n1177_n1297# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.5
.ends

.subckt isolated_switch_4 on off in vdd shunt out vss
XXM15 on m2_961_n2337# on on out on m2_961_n2337# m2_961_n2337# on m2_961_n2337# out
+ on vss out sky130_fd_pr__nfet_g5v0d10v5_F5JQJ7
XXM4 m2_961_n2337# out m2_961_n2337# off m2_961_n2337# out out off off off off off
+ off off off off off vdd m2_961_n2337# off out out m2_961_n2337# out m2_961_n2337#
+ out sky130_fd_pr__pfet_g5v0d10v5_AQSWZU
Xsky130_fd_pr__nfet_g5v0d10v5_F5JQJ7_0 on in on on m2_961_n2337# on in in on in m2_961_n2337#
+ on vss m2_961_n2337# sky130_fd_pr__nfet_g5v0d10v5_F5JQJ7
Xsky130_fd_pr__nfet_g5v0d10v5_EJGQJV_0 vss vss m2_961_n2337# shunt sky130_fd_pr__nfet_g5v0d10v5_EJGQJV
Xsky130_fd_pr__pfet_g5v0d10v5_AQSWZU_0 in m2_961_n2337# in off in m2_961_n2337# m2_961_n2337#
+ off off off off off off off off off off vdd in off m2_961_n2337# m2_961_n2337# in
+ m2_961_n2337# in m2_961_n2337# sky130_fd_pr__pfet_g5v0d10v5_AQSWZU
.ends

.subckt isolated_switch_xlarge on out in avdd off avss dvdd dvss
Xx2 on dvdd dvss avdd avdd x2/X avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xx3 off dvdd dvss avdd avdd x3/X avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xisolated_switch_4_0 x2/X isolated_switch_4_0/off in avdd x3/X out avss isolated_switch_4
Xsky130_fd_sc_hvl__diode_2_0 on dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_1 off dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_1_0 x2/X dvss dvss avdd avdd isolated_switch_4_0/off sky130_fd_sc_hvl__inv_1
.ends

.subckt switch_array_4 channel0_in_to_out[1] channel0_in_to_out[0] channel1_in_to_out[1]
+ channel1_in_to_out[0] channel2_in_to_out[1] channel2_in_to_out[0] channel3_in_to_out[1]
+ channel3_in_to_out[0] channel0_in channel0_out channel1_out channel2_in channel2_out
+ channel3_in channel3_out dvss avdd dvdd channel1_in avss
Xisolated_switch_xlarge_0[0|0] channel2_in_to_out[0] channel2_out channel2_in avdd
+ channel2_in_to_out[1] avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_0[1|0] channel3_in_to_out[0] channel3_out channel3_in avdd
+ channel3_in_to_out[1] avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_0[0|1] channel0_in_to_out[0] channel0_out channel0_in avdd
+ channel0_in_to_out[1] avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_0[1|1] channel1_in_to_out[0] channel1_out channel1_in avdd
+ channel1_in_to_out[1] avss dvdd dvss isolated_switch_xlarge
.ends

.subckt simple_switch_array_15 user_vinref vdda0 simplest_analog_switch_ena1v8_1[1]/on
+ comp_p simplest_analog_switch_ena1v8_1[0]/on isolated_switch_large_0[4]/off simplest_analog_switch_ena1v8_1[7]/on
+ simplest_analog_switch_ena1v8_1[5]/on comp_n left_vref isolated_switch_large_0[1]/off
+ isolated_switch_large_0[3]/on simplest_analog_switch_ena1v8_1[3]/on right_vref user_adc1
+ user_vbgsc dac1 user_adc0 user_vbgtc isolated_switch_large_0[0]/on dac0 vinref simplest_analog_switch_ena1v8_1[2]/on
+ tempsense isolated_switch_large_0[5]/off user_tempsense vbgsc vbgtc isolated_switch_large_0[4]/on
+ isolated_switch_large_0[2]/off simplest_analog_switch_ena1v8_1[8]/on isolated_switch_large_0[1]/on
+ user_dac1 user_dac0 simplest_analog_switch_ena1v8_1[6]/on ulpcomp_p user_left_vinref
+ simplest_analog_switch_ena1v8_1[4]/on ulpcomp_n isolated_switch_large_0[5]/on isolated_switch_large_0[3]/off
+ user_comp_p user_right_vinref user_ulpcomp_p user_comp_n isolated_switch_large_0[2]/on
+ isolated_switch_large_0[0]/off user_ulpcomp_n adc1 adc0 vccd0 voutref vssa0 vssd0
+ user_voutref
Xisolated_switch_large_0[0] vssa0 isolated_switch_large_0[0]/on vdda0 isolated_switch_large_0[0]/off
+ vccd0 user_ulpcomp_p ulpcomp_p vssd0 isolated_switch_large
Xisolated_switch_large_0[1] vssa0 isolated_switch_large_0[1]/on vdda0 isolated_switch_large_0[1]/off
+ vccd0 user_ulpcomp_n ulpcomp_n vssd0 isolated_switch_large
Xisolated_switch_large_0[2] vssa0 isolated_switch_large_0[2]/on vdda0 isolated_switch_large_0[2]/off
+ vccd0 user_comp_p comp_p vssd0 isolated_switch_large
Xisolated_switch_large_0[3] vssa0 isolated_switch_large_0[3]/on vdda0 isolated_switch_large_0[3]/off
+ vccd0 user_comp_n comp_n vssd0 isolated_switch_large
Xisolated_switch_large_0[4] vssa0 isolated_switch_large_0[4]/on vdda0 isolated_switch_large_0[4]/off
+ vccd0 user_adc1 adc1 vssd0 isolated_switch_large
Xisolated_switch_large_0[5] vssa0 isolated_switch_large_0[5]/on vdda0 isolated_switch_large_0[5]/off
+ vccd0 user_adc0 adc0 vssd0 isolated_switch_large
Xsimplest_analog_switch_ena1v8_1[0] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[0]/on
+ user_vbgsc vssd0 vbgsc simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[1]/on
+ user_vbgtc vssd0 vbgtc simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[2] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[2]/on
+ user_dac1 vssd0 dac1 simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[3] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[3]/on
+ user_dac0 vssd0 dac0 simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[4] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[4]/on
+ user_tempsense vssd0 tempsense simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[5] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[5]/on
+ user_right_vinref vssd0 right_vref simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[6] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[6]/on
+ user_left_vinref vssd0 left_vref simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[7] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[7]/on
+ user_vinref vssd0 vinref simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[8] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[8]/on
+ user_voutref vssd0 voutref simplest_analog_switch_ena1v8
.ends

.subckt simple_switch_array_8 simplest_analog_switch_ena1v8_1[3]/in simplest_analog_switch_ena1v8_1[2]/in
+ simplest_analog_switch_ena1v8_1[2]/on simplest_analog_switch_ena1v8_1[1]/on simplest_analog_switch_ena1v8_0[1]/in
+ simplest_analog_switch_ena1v8_0[0]/in simplest_analog_switch_ena1v8_0[3]/on simplest_analog_switch_ena1v8_0[0]/on
+ simplest_analog_switch_ena1v8_0[2]/on simplest_analog_switch_ena1v8_0[1]/on simplest_analog_switch_ena1v8_1[1]/in
+ simplest_analog_switch_ena1v8_0[3]/in simplest_analog_switch_ena1v8_1[0]/on simplest_analog_switch_ena1v8_1[0]/in
+ simplest_analog_switch_ena1v8_1[3]/on simplest_analog_switch_ena1v8_1[3]/dvdd simplest_analog_switch_ena1v8_1[3]/out
+ simplest_analog_switch_ena1v8_0[2]/in simplest_analog_switch_ena1v8_1[3]/avss simplest_analog_switch_ena1v8_0[3]/out
+ simplest_analog_switch_ena1v8_1[3]/avdd VSUBS
Xsimplest_analog_switch_ena1v8_0[0] simplest_analog_switch_ena1v8_1[3]/avdd simplest_analog_switch_ena1v8_1[3]/dvdd
+ simplest_analog_switch_ena1v8_1[3]/avss simplest_analog_switch_ena1v8_0[0]/on simplest_analog_switch_ena1v8_0[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[1] simplest_analog_switch_ena1v8_1[3]/avdd simplest_analog_switch_ena1v8_1[3]/dvdd
+ simplest_analog_switch_ena1v8_1[3]/avss simplest_analog_switch_ena1v8_0[1]/on simplest_analog_switch_ena1v8_0[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[2] simplest_analog_switch_ena1v8_1[3]/avdd simplest_analog_switch_ena1v8_1[3]/dvdd
+ simplest_analog_switch_ena1v8_1[3]/avss simplest_analog_switch_ena1v8_0[2]/on simplest_analog_switch_ena1v8_0[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[2]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[3] simplest_analog_switch_ena1v8_1[3]/avdd simplest_analog_switch_ena1v8_1[3]/dvdd
+ simplest_analog_switch_ena1v8_1[3]/avss simplest_analog_switch_ena1v8_0[3]/on simplest_analog_switch_ena1v8_0[3]/out
+ VSUBS simplest_analog_switch_ena1v8_0[3]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[0] simplest_analog_switch_ena1v8_1[3]/avdd simplest_analog_switch_ena1v8_1[3]/dvdd
+ simplest_analog_switch_ena1v8_1[3]/avss simplest_analog_switch_ena1v8_1[0]/on simplest_analog_switch_ena1v8_1[3]/out
+ VSUBS simplest_analog_switch_ena1v8_1[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1] simplest_analog_switch_ena1v8_1[3]/avdd simplest_analog_switch_ena1v8_1[3]/dvdd
+ simplest_analog_switch_ena1v8_1[3]/avss simplest_analog_switch_ena1v8_1[1]/on simplest_analog_switch_ena1v8_1[3]/out
+ VSUBS simplest_analog_switch_ena1v8_1[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[2] simplest_analog_switch_ena1v8_1[3]/avdd simplest_analog_switch_ena1v8_1[3]/dvdd
+ simplest_analog_switch_ena1v8_1[3]/avss simplest_analog_switch_ena1v8_1[2]/on simplest_analog_switch_ena1v8_1[3]/out
+ VSUBS simplest_analog_switch_ena1v8_1[2]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[3] simplest_analog_switch_ena1v8_1[3]/avdd simplest_analog_switch_ena1v8_1[3]/dvdd
+ simplest_analog_switch_ena1v8_1[3]/avss simplest_analog_switch_ena1v8_1[3]/on simplest_analog_switch_ena1v8_1[3]/out
+ VSUBS simplest_analog_switch_ena1v8_1[3]/in simplest_analog_switch_ena1v8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_9992MR__0 a_50_n136# a_n108_n136# a_n50_n162#
+ w_n144_n198#
X0 a_50_n136# a_n50_n162# a_n108_n136# w_n144_n198# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt poly_res_200ohm a_n414_974# a_n414_n76#
X0 a_n414_974# a_n414_n76# sky130_fd_pr__res_generic_po w=0.71 l=2.96
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0 a_n108_n34# a_n50_n122# a_50_n34# VSUBS
X0 a_50_n34# a_n50_n122# a_n108_n34# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.1885 pd=1.88 as=0.1885 ps=1.88 w=0.65 l=0.5
.ends

.subckt rheo_3v_cell_top m1_814_1199# w_318_n275# m1_545_847# m1_387_847# m1_824_799#
+ w_318_892# m1_290_1114# poly_res_200ohm_1/VSUBS m1_545_212# m1_663_847# m1_300_n125#
+ m4_97_801# m1_821_212# m4_97_1059# m1_814_483# poly_res_200ohm_0/a_n414_n76# m1_663_212#
+ m1_155_n223# m1_814_591# m1_814_n125# m1_290_591# m1_290_344#
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_545_847# m1_387_847# m1_290_1114# w_318_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_663_847# m1_814_1199# w_318_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_821_212# m1_663_212# m1_814_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xpoly_res_200ohm_0 m1_824_799# poly_res_200ohm_0/a_n414_n76# poly_res_200ohm
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# m1_300_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xpoly_res_200ohm_1 m1_824_799# m1_155_n223# poly_res_200ohm
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# m1_290_591# m1_545_847# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_663_847# m1_814_591# m1_824_799# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# m1_290_344# m1_545_212# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_663_212# m1_814_483# m1_821_212# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_9992MR a_50_n136# a_n108_n136# a_n50_n162# w_n144_n198#
X0 a_50_n136# a_n50_n162# a_n108_n136# w_n144_n198# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NHLDUY a_n108_n34# a_n50_n122# a_50_n34# VSUBS
X0 a_50_n34# a_n50_n122# a_n108_n34# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.1885 pd=1.88 as=0.1885 ps=1.88 w=0.65 l=0.5
.ends

.subckt rheo_3v_cell m1_814_1199# w_318_n275# m1_545_847# m1_387_847# m1_290_1114#
+ poly_res_200ohm_1/VSUBS m1_545_212# m1_663_847# m1_300_n125# m1_821_212# m1_824_799#
+ m1_814_483# poly_res_200ohm_1/a_n414_974# poly_res_200ohm_0/a_n414_n76# m1_663_212#
+ m1_155_n223# m1_814_591# w_316_892# m1_814_n125# m1_290_591# m1_290_344#
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_545_847# m1_387_847# m1_290_1114# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_663_847# m1_814_1199# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_821_212# m1_663_212# m1_814_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xpoly_res_200ohm_0 m1_824_799# poly_res_200ohm_0/a_n414_n76# poly_res_200ohm
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# m1_300_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xpoly_res_200ohm_1 poly_res_200ohm_1/a_n414_974# m1_155_n223# poly_res_200ohm
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# m1_290_591# m1_545_847# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_663_847# m1_814_591# m1_824_799# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# m1_290_344# m1_545_212# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_663_212# m1_814_483# m1_821_212# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
.ends

.subckt rheo_3v_column rheo_3v_cell_top_0/m4_97_1059# b3b b0_uq14 b0_uq3 b2b_uq1 dum1_out
+ b0_uq2 rheo_3v_cell_0[1]/w_316_892# b0b_uq14 b3 rheo_3v_cell_top_0/m1_290_591# b1_uq6
+ b0b_uq9 rheo_3v_cell_0[5]/w_316_892# b0_uq13 b0b_uq12 b1 rheo_3v_cell_0[6]/w_316_892#
+ b0b_uq8 dum0_in b0b_uq7 b2 b1_uq3 b0_uq0 b0b_uq6 b1_uq2 rheo_3v_cell_top_0/m1_290_1114#
+ b1_uq1 b1_uq5 b1_uq0 b3_uq0 b3b_uq0 b1_uq4 b0b_uq5 rheo_3v_cell_0[4]/w_316_892#
+ b0_uq5 m2_801_196# rheo_3v_cell_0[7]/w_316_892# b0b_uq0 b0b_uq13 b0_uq4 b0b_uq4
+ out_5 b0_uq11 b2b_uq0 out_4 b4 b0_uq10 rheo_3v_cell_0[3]/w_316_892# b2_uq2 b0b_uq3
+ b2_uq1 b0_uq12 m2_801_13759# res0_in b0b_uq1 b0b_uq2 b1b_uq3 b1b_uq4 b1b_uq6 b1b_uq2
+ b4b b1b_uq1 b2b_uq2 b1b_uq0 b1b_uq5 m2_791_1314# b2_uq0 b0b_uq11 rheo_3v_cell_0[2]/w_316_892#
+ b0_uq9 b0b b0_uq1 res1_out b0_uq8 rheo_3v_cell_top_0/m4_97_801# b0_uq6 b0b_uq10
+ m2_791_14877# b1b b0_uq7 b0 b2b VSUBS
Xrheo_3v_cell_top_0 b0_uq14 rheo_3v_cell_0[7]/w_316_892# out_4 out_5 res1_in m2_801_13759#
+ rheo_3v_cell_top_0/m1_290_1114# VSUBS out0_0_3 out1_0_0 b0b_uq13 rheo_3v_cell_top_0/m4_97_801#
+ out1_1_0 rheo_3v_cell_top_0/m4_97_1059# b1_uq6 rheo_3v_cell_0[7]/m1_824_799# out1_0_0
+ rheo_3v_cell_top_0/m1_155_n223# b0b_uq14 b1b_uq6 rheo_3v_cell_top_0/m1_290_591#
+ b0_uq13 rheo_3v_cell_top
Xrheo_3v_cell_0[0] m2_791_1314# m2_801_196# m2_328_1119# m2_328_1119# m2_791_1314#
+ VSUBS m2_449_485# m2_328_1119# m2_801_196# m2_449_485# res1_out VSUBS res0_in dum1_out
+ m2_449_485# dum0_in VSUBS m2_791_1314# m2_801_196# VSUBS VSUBS rheo_3v_cell
Xrheo_3v_cell_0[1] b0b m2_791_1314# out0_0_0 out0_1_0 b1b_uq0 VSUBS out0_0_0 out1_0_3
+ b0_uq0 out_3 rheo_3v_cell_0[1]/m1_824_799# b4b rheo_3v_cell_0[2]/m1_155_n223# res1_out
+ out_4 res0_in b0 rheo_3v_cell_0[1]/w_316_892# b4 b1_uq0 b0b_uq0 rheo_3v_cell
Xrheo_3v_cell_0[2] b0_uq2 rheo_3v_cell_0[1]/w_316_892# out0_2 out0_1_0 b2b_uq0 VSUBS
+ out0_0_0 out1_0_3 b0b_uq1 out1_1_1 rheo_3v_cell_0[2]/m1_824_799# b1b rheo_3v_cell_0[3]/m1_155_n223#
+ rheo_3v_cell_0[1]/m1_824_799# out1_0_3 rheo_3v_cell_0[2]/m1_155_n223# b0b_uq2 rheo_3v_cell_0[2]/w_316_892#
+ b1 b2_uq0 b0_uq1 rheo_3v_cell
Xrheo_3v_cell_0[3] b0b_uq4 rheo_3v_cell_0[2]/w_316_892# out0_0_1 out0_1_0 b1_uq1 VSUBS
+ out0_0_1 out1_0_2 b0_uq3 out1_1_1 rheo_3v_cell_0[3]/m1_824_799# b2b rheo_3v_cell_0[4]/m1_155_n223#
+ rheo_3v_cell_0[2]/m1_824_799# out1_2 rheo_3v_cell_0[3]/m1_155_n223# b0_uq4 rheo_3v_cell_0[3]/w_316_892#
+ b2 b1b_uq1 b0b_uq3 rheo_3v_cell
Xrheo_3v_cell_0[4] b0_uq6 rheo_3v_cell_0[3]/w_316_892# out_3 out0_2 b3b_uq0 VSUBS
+ out0_0_1 out1_0_2 b0b_uq5 out1_1_1 rheo_3v_cell_0[4]/m1_824_799# b1_uq2 rheo_3v_cell_0[5]/m1_155_n223#
+ rheo_3v_cell_0[3]/m1_824_799# out1_0_2 rheo_3v_cell_0[4]/m1_155_n223# b0b_uq6 rheo_3v_cell_0[4]/w_316_892#
+ b1b_uq2 b3_uq0 b0_uq5 rheo_3v_cell
Xrheo_3v_cell_0[5] b0b_uq8 rheo_3v_cell_0[4]/w_316_892# out0_0_2 out0_1_1 b1b_uq3
+ VSUBS out0_0_2 out1_0_1 b0_uq7 out1_2 rheo_3v_cell_0[5]/m1_824_799# b3b rheo_3v_cell_0[6]/m1_155_n223#
+ rheo_3v_cell_0[4]/m1_824_799# out_3 rheo_3v_cell_0[5]/m1_155_n223# b0_uq8 rheo_3v_cell_0[5]/w_316_892#
+ b3 b1_uq3 b0b_uq7 rheo_3v_cell
Xrheo_3v_cell_0[6] b0_uq10 rheo_3v_cell_0[5]/w_316_892# out0_2 out0_1_1 b2_uq1 VSUBS
+ out0_0_2 out1_0_1 b0b_uq9 out1_1_0 rheo_3v_cell_0[6]/m1_824_799# b1b_uq4 rheo_3v_cell_0[7]/m1_155_n223#
+ rheo_3v_cell_0[5]/m1_824_799# out1_0_1 rheo_3v_cell_0[6]/m1_155_n223# b0b_uq10 rheo_3v_cell_0[6]/w_316_892#
+ b1_uq4 b2b_uq1 b0_uq9 rheo_3v_cell
Xrheo_3v_cell_0[7] b0b_uq12 rheo_3v_cell_0[6]/w_316_892# out0_0_3 out0_1_1 b1_uq5
+ VSUBS out0_0_3 out1_0_0 b0_uq11 out1_1_0 rheo_3v_cell_0[7]/m1_824_799# b2_uq2 rheo_3v_cell_top_0/m1_155_n223#
+ rheo_3v_cell_0[6]/m1_824_799# out1_2 rheo_3v_cell_0[7]/m1_155_n223# b0_uq12 rheo_3v_cell_0[7]/w_316_892#
+ b2b_uq2 b1b_uq5 b0b_uq11 rheo_3v_cell
Xrheo_3v_cell_1 m2_791_14877# m2_801_13759# m2_330_14682# m2_330_14682# m2_791_14877#
+ VSUBS m2_449_14048# m2_330_14682# m2_801_13759# m2_449_14048# dum0_out VSUBS dum0_out
+ res1_in m2_449_14048# res1_in VSUBS m2_791_14877# m2_801_13759# VSUBS VSUBS rheo_3v_cell
.ends

.subckt rheo_3v_cell_odd m1_814_1199# w_318_n275# m1_545_847# m1_387_847# m1_290_1114#
+ poly_res_200ohm_1/VSUBS m1_545_212# m1_663_847# m1_300_n125# m1_821_212# m1_824_799#
+ m1_814_483# poly_res_200ohm_1/a_n414_974# poly_res_200ohm_0/a_n414_n76# m1_663_212#
+ m1_155_n223# m1_814_591# w_316_892# m1_814_n125# m1_290_591# m1_290_344#
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_545_847# m1_387_847# m1_290_1114# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_663_847# m1_814_1199# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_821_212# m1_663_212# m1_814_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xpoly_res_200ohm_0 m1_824_799# poly_res_200ohm_0/a_n414_n76# poly_res_200ohm
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# m1_300_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xpoly_res_200ohm_1 poly_res_200ohm_1/a_n414_974# m1_155_n223# poly_res_200ohm
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# m1_290_591# m1_545_847# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_663_847# m1_814_591# m1_824_799# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# m1_290_344# m1_545_212# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_663_212# m1_814_483# m1_821_212# poly_res_200ohm_1/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
.ends

.subckt rheo_3v_column_odd rheo_3v_cell_top_0/m4_97_1059# m3_31_13582# res_in0 b0_uq14
+ b2b_uq2 b0_uq12 b0_uq6 rheo_3v_cell_0[1]/w_316_892# b0b_uq14 b1_uq6 rheo_3v_cell_0[0]/w_316_892#
+ b0_uq1 b0_uq13 b0b_uq12 b1 in_5 b0b_uq11 b3 b0b_uq10 b0_uq3 b3b b1_uq1 m3_30_13212#
+ b0_uq2 b0b_uq3 b2b_uq1 b0_uq0 b0b_uq9 rheo_3v_cell_0[4]/w_316_892# b0b_uq2 rheo_3v_cell_odd_0/w_316_892#
+ rheo_3v_cell_0[5]/w_316_892# b0b_uq1 b0b_uq13 b0b_uq8 b3b_uq0 b1_uq2 b4 b2 out_5
+ b1_uq3 dum_in0 res_out1 rheo_3v_cell_0[3]/w_316_892# b2_uq2 b0b_uq7 b1_uq5 b4b out4
+ b1b_uq5 b2_uq1 b1_uq4 m2_801_196# m2_791_14877# m2_801_13759# b1b_uq4 b0b_uq6 b0b_uq5
+ b0 b2_uq0 b1b_uq3 b1b_uq6 b1b_uq2 b0b_uq4 b1b_uq1 b1b_uq0 b0_uq11 b2b_uq0 b3_uq0
+ b1_uq0 rheo_3v_cell_0[2]/w_316_892# b0_uq9 dum_out1 b0_uq5 b0b b0b_uq0 b0_uq8 rheo_3v_cell_top_0/m4_97_801#
+ b0_uq10 m2_791_1314# b1b VSUBS b0_uq7 b0_uq4 b2b
Xrheo_3v_cell_2 m2_791_14877# m2_801_13759# m2_331_14682# m2_331_14682# m2_791_14877#
+ VSUBS m2_458_14048# m2_331_14682# m2_801_13759# m2_458_14048# dum_out0 VSUBS dum_out0
+ res_in1 m2_458_14048# res_in1 VSUBS m2_791_14877# m2_801_13759# VSUBS VSUBS rheo_3v_cell
Xrheo_3v_cell_odd_0 b0b m2_791_1314# out0_0_0 out0_1_0 b1b_uq0 VSUBS out0_0_0 out1_0_3
+ b0_uq0 out_3 rheo_3v_cell_odd_0/m1_824_799# b4 rheo_3v_cell_0[0]/m1_155_n223# res_out1
+ out4 res_in0 b0 rheo_3v_cell_odd_0/w_316_892# b4b b1_uq0 b0b_uq0 rheo_3v_cell_odd
Xrheo_3v_cell_top_0 b0_uq14 rheo_3v_cell_0[5]/w_316_892# in_5 out_5 res_in1 m2_801_13759#
+ m3_31_13582# VSUBS out0_0_3 out1_0_0 b0b_uq13 rheo_3v_cell_top_0/m4_97_801# out1_1_0
+ rheo_3v_cell_top_0/m4_97_1059# b1_uq6 rheo_3v_cell_0[5]/m1_824_799# out1_0_0 rheo_3v_cell_top_0/m1_155_n223#
+ b0b_uq14 b1b_uq6 m3_30_13212# b0_uq13 rheo_3v_cell_top
Xrheo_3v_cell_0[0] b0_uq2 rheo_3v_cell_odd_0/w_316_892# out0_2 out0_1_0 b2b_uq0 VSUBS
+ out0_0_0 out1_0_3 b0b_uq1 out1_1_1 rheo_3v_cell_0[0]/m1_824_799# b1b rheo_3v_cell_0[1]/m1_155_n223#
+ rheo_3v_cell_odd_0/m1_824_799# out1_0_3 rheo_3v_cell_0[0]/m1_155_n223# b0b_uq2 rheo_3v_cell_0[0]/w_316_892#
+ b1 b2_uq0 b0_uq1 rheo_3v_cell
Xrheo_3v_cell_0[1] b0b_uq4 rheo_3v_cell_0[0]/w_316_892# out0_0_1 out0_1_0 b1_uq1 VSUBS
+ out0_0_1 out1_0_2 b0_uq3 out1_1_1 rheo_3v_cell_0[1]/m1_824_799# b2b rheo_3v_cell_0[2]/m1_155_n223#
+ rheo_3v_cell_0[0]/m1_824_799# out1_2 rheo_3v_cell_0[1]/m1_155_n223# b0_uq4 rheo_3v_cell_0[1]/w_316_892#
+ b2 b1b_uq1 b0b_uq3 rheo_3v_cell
Xrheo_3v_cell_0[2] b0_uq6 rheo_3v_cell_0[1]/w_316_892# out_3 out0_2 b3b_uq0 VSUBS
+ out0_0_1 out1_0_2 b0b_uq5 out1_1_1 rheo_3v_cell_0[2]/m1_824_799# b1_uq2 rheo_3v_cell_0[3]/m1_155_n223#
+ rheo_3v_cell_0[1]/m1_824_799# out1_0_2 rheo_3v_cell_0[2]/m1_155_n223# b0b_uq6 rheo_3v_cell_0[2]/w_316_892#
+ b1b_uq2 b3_uq0 b0_uq5 rheo_3v_cell
Xrheo_3v_cell_0[3] b0b_uq8 rheo_3v_cell_0[2]/w_316_892# out0_0_2 m3_296_8710# b1b_uq3
+ VSUBS out0_0_2 out1_0_1 b0_uq7 out1_2 rheo_3v_cell_0[3]/m1_824_799# b3b rheo_3v_cell_0[4]/m1_155_n223#
+ rheo_3v_cell_0[2]/m1_824_799# out_3 rheo_3v_cell_0[3]/m1_155_n223# b0_uq8 rheo_3v_cell_0[3]/w_316_892#
+ b3 b1_uq3 b0b_uq7 rheo_3v_cell
Xrheo_3v_cell_0[4] b0_uq10 rheo_3v_cell_0[3]/w_316_892# out0_2 m3_296_8710# b2_uq1
+ VSUBS out0_0_2 out1_0_1 b0b_uq9 out1_1_0 rheo_3v_cell_0[4]/m1_824_799# b1b_uq4 rheo_3v_cell_0[5]/m1_155_n223#
+ rheo_3v_cell_0[3]/m1_824_799# out1_0_1 rheo_3v_cell_0[4]/m1_155_n223# b0b_uq10 rheo_3v_cell_0[4]/w_316_892#
+ b1_uq4 b2b_uq1 b0_uq9 rheo_3v_cell
Xrheo_3v_cell_0[5] b0b_uq12 rheo_3v_cell_0[4]/w_316_892# out0_0_3 m3_296_8710# b1_uq5
+ VSUBS out0_0_3 out1_0_0 b0_uq11 out1_1_0 rheo_3v_cell_0[5]/m1_824_799# b2_uq2 rheo_3v_cell_top_0/m1_155_n223#
+ rheo_3v_cell_0[4]/m1_824_799# out1_2 rheo_3v_cell_0[5]/m1_155_n223# b0_uq12 rheo_3v_cell_0[5]/w_316_892#
+ b2b_uq2 b1b_uq5 b0b_uq11 rheo_3v_cell
Xrheo_3v_cell_1 m2_791_1314# m2_801_196# m2_329_1119# m2_329_1119# m2_791_1314# VSUBS
+ m2_457_485# m2_329_1119# m2_801_196# m2_457_485# res_out1 VSUBS res_in0 dum_out1
+ m2_457_485# dum_in0 VSUBS m2_791_1314# m2_801_196# VSUBS VSUBS rheo_3v_cell
.ends

.subckt rheo_3v_cell_dummy m4_99_18# w_318_n275# m4_99_276# m4_99_801# poly_res_200ohm_1/VSUBS
+ m4_99_930# m1_824_799# poly_res_200ohm_1/a_n414_974# m4_99_405# m4_99_1059# poly_res_200ohm_0/a_n414_n76#
+ m4_99_672# m1_155_n223# w_316_892# m4_99_147#
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_387_847# m1_387_847# w_316_892# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_387_847# w_316_892# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_545_212# m1_545_212# w_318_n275# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xpoly_res_200ohm_0 m1_824_799# poly_res_200ohm_0/a_n414_n76# poly_res_200ohm
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# w_318_n275# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR
Xpoly_res_200ohm_1 poly_res_200ohm_1/a_n414_974# m1_155_n223# poly_res_200ohm
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# poly_res_200ohm_1/VSUBS m1_387_847#
+ poly_res_200ohm_1/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_387_847# poly_res_200ohm_1/VSUBS m1_824_799#
+ poly_res_200ohm_1/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# poly_res_200ohm_1/VSUBS m1_545_212#
+ poly_res_200ohm_1/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_545_212# poly_res_200ohm_1/VSUBS m1_545_212#
+ poly_res_200ohm_1/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY
.ends

.subckt rheo_3v_column_dummy rheo_3v_cell_dummy_0[7]/m4_99_930# rheo_3v_cell_dummy_0[7]/m4_99_1059#
+ rheo_3v_cell_dummy_0[2]/m4_99_1059# rheo_3v_cell_dummy_0[8]/m4_99_18# rheo_3v_cell_dummy_0[8]/m4_99_930#
+ rheo_3v_cell_dummy_0[0]/m4_99_405# rheo_3v_cell_dummy_0[9]/m4_99_930# rheo_3v_cell_dummy_0[1]/m4_99_405#
+ rheo_3v_cell_dummy_0[2]/m4_99_405# rheo_3v_cell_dummy_0[0]/m4_99_672# rheo_3v_cell_dummy_0[9]/m4_99_18#
+ rheo_3v_cell_dummy_0[1]/m4_99_672# rheo_3v_cell_dummy_0[3]/m4_99_405# rheo_3v_cell_dummy_0[2]/m4_99_672#
+ rheo_3v_cell_dummy_0[4]/m4_99_405# rheo_3v_cell_dummy_0[5]/m4_99_405# rheo_3v_cell_dummy_0[3]/m4_99_672#
+ rheo_3v_cell_dummy_0[6]/m4_99_405# rheo_3v_cell_dummy_0[4]/m4_99_672# rheo_3v_cell_dummy_0[3]/w_316_892#
+ rheo_3v_cell_dummy_0[5]/m4_99_672# rheo_3v_cell_dummy_0[7]/m4_99_405# rheo_3v_cell_dummy_0[6]/m4_99_1059#
+ rheo_3v_cell_dummy_0[1]/m4_99_1059# rheo_3v_cell_dummy_0[8]/m4_99_405# rheo_3v_cell_dummy_0[6]/m4_99_672#
+ rheo_3v_cell_dummy_0[7]/m4_99_672# rheo_3v_cell_dummy_0[9]/m4_99_405# rheo_3v_cell_dummy_0[2]/w_316_892#
+ rheo_3v_cell_dummy_0[8]/m4_99_672# rheo_3v_cell_dummy_0[0]/m4_99_18# rheo_3v_cell_dummy_0[0]/m4_99_147#
+ rheo_3v_cell_dummy_0[7]/w_316_892# rheo_3v_cell_dummy_0[9]/m4_99_672# rheo_3v_cell_dummy_0[8]/w_316_892#
+ rheo_3v_cell_dummy_0[1]/m4_99_147# rheo_3v_cell_dummy_0[9]/w_316_892# rheo_3v_cell_dummy_0[2]/m4_99_147#
+ rheo_3v_cell_dummy_0[3]/m4_99_147# rheo_3v_cell_dummy_0[1]/m4_99_18# rheo_3v_cell_dummy_0[4]/m4_99_147#
+ rheo_3v_cell_dummy_0[5]/m4_99_147# rheo_3v_cell_dummy_0[5]/m4_99_1059# rheo_3v_cell_dummy_0[0]/m4_99_1059#
+ rheo_3v_cell_dummy_0[6]/m4_99_147# rheo_3v_cell_dummy_0[6]/w_316_892# rheo_3v_cell_dummy_0[7]/m4_99_147#
+ rheo_3v_cell_dummy_0[1]/w_316_892# rheo_3v_cell_dummy_0[2]/m4_99_18# rheo_3v_cell_dummy_0[8]/m4_99_147#
+ rheo_3v_cell_dummy_0[9]/m4_99_147# rheo_3v_cell_dummy_0[3]/m4_99_18# rheo_3v_cell_dummy_0[0]/m4_99_276#
+ rheo_3v_cell_dummy_0[0]/m4_99_801# rheo_3v_cell_dummy_0[1]/m4_99_276# rheo_3v_cell_dummy_0[9]/m4_99_1059#
+ rheo_3v_cell_dummy_0[1]/m4_99_801# rheo_3v_cell_dummy_0[4]/m4_99_1059# rheo_3v_cell_dummy_0[2]/m4_99_276#
+ rheo_3v_cell_dummy_0[2]/m4_99_801# rheo_3v_cell_dummy_0[3]/m4_99_276# rheo_3v_cell_dummy_0[3]/m4_99_801#
+ rheo_3v_cell_dummy_0[5]/w_316_892# rheo_3v_cell_dummy_0[4]/m4_99_18# rheo_3v_cell_dummy_0[4]/m4_99_276#
+ rheo_3v_cell_dummy_0[0]/w_316_892# rheo_3v_cell_dummy_0[4]/m4_99_801# rheo_3v_cell_dummy_0[5]/m4_99_276#
+ rheo_3v_cell_dummy_0[5]/m4_99_801# rheo_3v_cell_dummy_0[6]/m4_99_276# rheo_3v_cell_dummy_0[6]/m4_99_801#
+ rheo_3v_cell_dummy_0[7]/m4_99_276# rheo_3v_cell_dummy_0[7]/m4_99_801# rheo_3v_cell_dummy_0[8]/m4_99_276#
+ rheo_3v_cell_dummy_0[5]/m4_99_18# rheo_3v_cell_dummy_0[8]/m4_99_801# rheo_3v_cell_dummy_0[9]/m4_99_276#
+ rheo_3v_cell_dummy_0[9]/m4_99_801# rheo_3v_cell_dummy_0[8]/m4_99_1059# rheo_3v_cell_dummy_0[3]/m4_99_1059#
+ rheo_3v_cell_dummy_0[6]/m4_99_18# rheo_3v_cell_dummy_0[0]/m4_99_930# rheo_3v_cell_dummy_0[4]/w_316_892#
+ rheo_3v_cell_dummy_0[0]/w_318_n275# rheo_3v_cell_dummy_0[1]/m4_99_930# rheo_3v_cell_dummy_0[2]/m4_99_930#
+ m1_988_1608# rheo_3v_cell_dummy_0[3]/m4_99_930# rheo_3v_cell_dummy_0[7]/m4_99_18#
+ m1_n18_1607# rheo_3v_cell_dummy_0[4]/m4_99_930# m1_938_45# rheo_3v_cell_dummy_0[5]/m4_99_930#
+ rheo_3v_cell_dummy_0[6]/m4_99_930# m1_n18_45# VSUBS
Xrheo_3v_cell_dummy_0[0] rheo_3v_cell_dummy_0[0]/m4_99_18# rheo_3v_cell_dummy_0[0]/w_318_n275#
+ rheo_3v_cell_dummy_0[0]/m4_99_276# rheo_3v_cell_dummy_0[0]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[0]/m4_99_930#
+ m1_988_1608# m1_n18_1607# rheo_3v_cell_dummy_0[0]/m4_99_405# rheo_3v_cell_dummy_0[0]/m4_99_1059#
+ m1_938_45# rheo_3v_cell_dummy_0[0]/m4_99_672# m1_n18_45# rheo_3v_cell_dummy_0[0]/w_316_892#
+ rheo_3v_cell_dummy_0[0]/m4_99_147# rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[1] rheo_3v_cell_dummy_0[1]/m4_99_18# rheo_3v_cell_dummy_0[0]/w_316_892#
+ rheo_3v_cell_dummy_0[1]/m4_99_276# rheo_3v_cell_dummy_0[1]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[1]/m4_99_930#
+ rheo_3v_cell_dummy_0[1]/m1_824_799# rheo_3v_cell_dummy_0[2]/m1_155_n223# rheo_3v_cell_dummy_0[1]/m4_99_405#
+ rheo_3v_cell_dummy_0[1]/m4_99_1059# m1_988_1608# rheo_3v_cell_dummy_0[1]/m4_99_672#
+ m1_n18_1607# rheo_3v_cell_dummy_0[1]/w_316_892# rheo_3v_cell_dummy_0[1]/m4_99_147#
+ rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[2] rheo_3v_cell_dummy_0[2]/m4_99_18# rheo_3v_cell_dummy_0[1]/w_316_892#
+ rheo_3v_cell_dummy_0[2]/m4_99_276# rheo_3v_cell_dummy_0[2]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[2]/m4_99_930#
+ rheo_3v_cell_dummy_0[2]/m1_824_799# rheo_3v_cell_dummy_0[3]/m1_155_n223# rheo_3v_cell_dummy_0[2]/m4_99_405#
+ rheo_3v_cell_dummy_0[2]/m4_99_1059# rheo_3v_cell_dummy_0[1]/m1_824_799# rheo_3v_cell_dummy_0[2]/m4_99_672#
+ rheo_3v_cell_dummy_0[2]/m1_155_n223# rheo_3v_cell_dummy_0[2]/w_316_892# rheo_3v_cell_dummy_0[2]/m4_99_147#
+ rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[3] rheo_3v_cell_dummy_0[3]/m4_99_18# rheo_3v_cell_dummy_0[2]/w_316_892#
+ rheo_3v_cell_dummy_0[3]/m4_99_276# rheo_3v_cell_dummy_0[3]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[3]/m4_99_930#
+ rheo_3v_cell_dummy_0[3]/m1_824_799# rheo_3v_cell_dummy_0[4]/m1_155_n223# rheo_3v_cell_dummy_0[3]/m4_99_405#
+ rheo_3v_cell_dummy_0[3]/m4_99_1059# rheo_3v_cell_dummy_0[2]/m1_824_799# rheo_3v_cell_dummy_0[3]/m4_99_672#
+ rheo_3v_cell_dummy_0[3]/m1_155_n223# rheo_3v_cell_dummy_0[3]/w_316_892# rheo_3v_cell_dummy_0[3]/m4_99_147#
+ rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[4] rheo_3v_cell_dummy_0[4]/m4_99_18# rheo_3v_cell_dummy_0[3]/w_316_892#
+ rheo_3v_cell_dummy_0[4]/m4_99_276# rheo_3v_cell_dummy_0[4]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[4]/m4_99_930#
+ rheo_3v_cell_dummy_0[4]/m1_824_799# rheo_3v_cell_dummy_0[5]/m1_155_n223# rheo_3v_cell_dummy_0[4]/m4_99_405#
+ rheo_3v_cell_dummy_0[4]/m4_99_1059# rheo_3v_cell_dummy_0[3]/m1_824_799# rheo_3v_cell_dummy_0[4]/m4_99_672#
+ rheo_3v_cell_dummy_0[4]/m1_155_n223# rheo_3v_cell_dummy_0[4]/w_316_892# rheo_3v_cell_dummy_0[4]/m4_99_147#
+ rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[5] rheo_3v_cell_dummy_0[5]/m4_99_18# rheo_3v_cell_dummy_0[4]/w_316_892#
+ rheo_3v_cell_dummy_0[5]/m4_99_276# rheo_3v_cell_dummy_0[5]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[5]/m4_99_930#
+ rheo_3v_cell_dummy_0[5]/m1_824_799# rheo_3v_cell_dummy_0[6]/m1_155_n223# rheo_3v_cell_dummy_0[5]/m4_99_405#
+ rheo_3v_cell_dummy_0[5]/m4_99_1059# rheo_3v_cell_dummy_0[4]/m1_824_799# rheo_3v_cell_dummy_0[5]/m4_99_672#
+ rheo_3v_cell_dummy_0[5]/m1_155_n223# rheo_3v_cell_dummy_0[5]/w_316_892# rheo_3v_cell_dummy_0[5]/m4_99_147#
+ rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[6] rheo_3v_cell_dummy_0[6]/m4_99_18# rheo_3v_cell_dummy_0[5]/w_316_892#
+ rheo_3v_cell_dummy_0[6]/m4_99_276# rheo_3v_cell_dummy_0[6]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[6]/m4_99_930#
+ rheo_3v_cell_dummy_0[6]/m1_824_799# rheo_3v_cell_dummy_0[7]/m1_155_n223# rheo_3v_cell_dummy_0[6]/m4_99_405#
+ rheo_3v_cell_dummy_0[6]/m4_99_1059# rheo_3v_cell_dummy_0[5]/m1_824_799# rheo_3v_cell_dummy_0[6]/m4_99_672#
+ rheo_3v_cell_dummy_0[6]/m1_155_n223# rheo_3v_cell_dummy_0[6]/w_316_892# rheo_3v_cell_dummy_0[6]/m4_99_147#
+ rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[7] rheo_3v_cell_dummy_0[7]/m4_99_18# rheo_3v_cell_dummy_0[6]/w_316_892#
+ rheo_3v_cell_dummy_0[7]/m4_99_276# rheo_3v_cell_dummy_0[7]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[7]/m4_99_930#
+ rheo_3v_cell_dummy_0[7]/m1_824_799# rheo_3v_cell_dummy_0[8]/m1_155_n223# rheo_3v_cell_dummy_0[7]/m4_99_405#
+ rheo_3v_cell_dummy_0[7]/m4_99_1059# rheo_3v_cell_dummy_0[6]/m1_824_799# rheo_3v_cell_dummy_0[7]/m4_99_672#
+ rheo_3v_cell_dummy_0[7]/m1_155_n223# rheo_3v_cell_dummy_0[7]/w_316_892# rheo_3v_cell_dummy_0[7]/m4_99_147#
+ rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[8] rheo_3v_cell_dummy_0[8]/m4_99_18# rheo_3v_cell_dummy_0[7]/w_316_892#
+ rheo_3v_cell_dummy_0[8]/m4_99_276# rheo_3v_cell_dummy_0[8]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[8]/m4_99_930#
+ m1_36_13186# m1_36_13186# rheo_3v_cell_dummy_0[8]/m4_99_405# rheo_3v_cell_dummy_0[8]/m4_99_1059#
+ rheo_3v_cell_dummy_0[7]/m1_824_799# rheo_3v_cell_dummy_0[8]/m4_99_672# rheo_3v_cell_dummy_0[8]/m1_155_n223#
+ rheo_3v_cell_dummy_0[8]/w_316_892# rheo_3v_cell_dummy_0[8]/m4_99_147# rheo_3v_cell_dummy
Xrheo_3v_cell_dummy_0[9] rheo_3v_cell_dummy_0[9]/m4_99_18# rheo_3v_cell_dummy_0[8]/w_316_892#
+ rheo_3v_cell_dummy_0[9]/m4_99_276# rheo_3v_cell_dummy_0[9]/m4_99_801# VSUBS rheo_3v_cell_dummy_0[9]/m4_99_930#
+ m1_28_15111# m1_28_15111# rheo_3v_cell_dummy_0[9]/m4_99_405# rheo_3v_cell_dummy_0[9]/m4_99_1059#
+ m1_36_13186# rheo_3v_cell_dummy_0[9]/m4_99_672# m1_36_13186# rheo_3v_cell_dummy_0[9]/w_316_892#
+ rheo_3v_cell_dummy_0[9]/m4_99_147# rheo_3v_cell_dummy
.ends

.subckt sky130_fd_sc_hvl__inv_8 A VGND VNB VPB VPWR Y
X0 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.1575 pd=1.17 as=0.105 ps=1.03 w=0.75 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.20625 pd=2.05 as=0.105 ps=1.03 w=0.75 l=0.5
X3 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X4 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X5 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X6 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X7 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.1575 ps=1.17 w=0.75 l=0.5
X8 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X9 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X10 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X11 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X12 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X13 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X14 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X15 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
.ends

.subckt sky130_fd_sc_hvl__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X1 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X3 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.4275 ps=3.57 w=1.5 l=0.5
X4 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X5 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X7 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_4AXGXB a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt rheo_level_shifter dvdd avdd bitb_out bit_out bit_in agnd
Xsky130_fd_sc_hvl__inv_8_1 bitb_out agnd agnd avdd avdd bit_out sky130_fd_sc_hvl__inv_8
Xsky130_fd_sc_hvl__inv_4_0 sky130_fd_sc_hvl__inv_4_0/A agnd agnd avdd avdd sky130_fd_sc_hvl__inv_8_0/A
+ sky130_fd_sc_hvl__inv_4
Xsky130_fd_sc_hvl__inv_2_0 sky130_fd_sc_hvl__inv_2_0/A agnd agnd avdd avdd sky130_fd_sc_hvl__inv_4_0/A
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 bit_in dvdd agnd avdd avdd sky130_fd_sc_hvl__inv_2_0/A
+ avdd agnd agnd sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_pr__diode_pw2nd_05v5_4AXGXB_0 agnd bit_in sky130_fd_pr__diode_pw2nd_05v5_4AXGXB
Xsky130_fd_sc_hvl__inv_8_0 sky130_fd_sc_hvl__inv_8_0/A agnd agnd avdd avdd bitb_out
+ sky130_fd_sc_hvl__inv_8
.ends

.subckt rheo_level_shifter_array rheo_level_shifter_0[0]/bit_in rheo_level_shifter_0[3]/bit_out
+ rheo_level_shifter_0[3]/bitb_out rheo_level_shifter_0[4]/bit_in rheo_level_shifter_0[0]/bit_out
+ rheo_level_shifter_0[4]/bitb_out rheo_level_shifter_0[7]/bit_out rheo_level_shifter_0[1]/bit_in
+ rheo_level_shifter_0[0]/bitb_out rheo_level_shifter_0[5]/bit_in rheo_level_shifter_0[4]/bit_out
+ rheo_level_shifter_0[7]/bitb_out rheo_level_shifter_0[1]/bit_out rheo_level_shifter_0[5]/bitb_out
+ rheo_level_shifter_0[1]/bitb_out rheo_level_shifter_0[6]/bit_in rheo_level_shifter_0[2]/bit_in
+ rheo_level_shifter_0[5]/bit_out rheo_level_shifter_0[6]/bitb_out rheo_level_shifter_0[2]/bit_out
+ rheo_level_shifter_0[2]/bitb_out rheo_level_shifter_0[3]/bit_in rheo_level_shifter_0[7]/bit_in
+ rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd rheo_level_shifter_0[6]/bit_out
+ VSUBS
Xrheo_level_shifter_0[0] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[0]/bitb_out rheo_level_shifter_0[0]/bit_out rheo_level_shifter_0[0]/bit_in
+ VSUBS rheo_level_shifter
Xrheo_level_shifter_0[1] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[1]/bitb_out rheo_level_shifter_0[1]/bit_out rheo_level_shifter_0[1]/bit_in
+ VSUBS rheo_level_shifter
Xrheo_level_shifter_0[2] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[2]/bitb_out rheo_level_shifter_0[2]/bit_out rheo_level_shifter_0[2]/bit_in
+ VSUBS rheo_level_shifter
Xrheo_level_shifter_0[3] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[3]/bitb_out rheo_level_shifter_0[3]/bit_out rheo_level_shifter_0[3]/bit_in
+ VSUBS rheo_level_shifter
Xrheo_level_shifter_0[4] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[4]/bitb_out rheo_level_shifter_0[4]/bit_out rheo_level_shifter_0[4]/bit_in
+ VSUBS rheo_level_shifter
Xrheo_level_shifter_0[5] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[5]/bitb_out rheo_level_shifter_0[5]/bit_out rheo_level_shifter_0[5]/bit_in
+ VSUBS rheo_level_shifter
Xrheo_level_shifter_0[6] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[6]/bitb_out rheo_level_shifter_0[6]/bit_out rheo_level_shifter_0[6]/bit_in
+ VSUBS rheo_level_shifter
Xrheo_level_shifter_0[7] rheo_level_shifter_0[7]/dvdd rheo_level_shifter_0[7]/avdd
+ rheo_level_shifter_0[7]/bitb_out rheo_level_shifter_0[7]/bit_out rheo_level_shifter_0[7]/bit_in
+ VSUBS rheo_level_shifter
.ends

.subckt sky130_ef_ip__rheostat_8bit b0 b1 b2 b3 b4 b5 b6 b7 out vdd dvdd Vhigh vss
+ Vlow dvss
Xrheo_3v_column_0 b5a b3a b0b b0b b2a rheo_3v_column_0/dum1_out b0b vdd b0a b3b b5b
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_0/dum0_in b0a b2b b1b b0b b0a b1b
+ b5a b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_1/out_5
+ b0b b2a rheo_3v_column_0/out_4 b4a b0b vdd b2b b0a b2b b0b vdd Vhigh b0a b0a b1a
+ b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_0/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_1 b5a b3a b0b b0b b2a rheo_3v_column_1/dum1_out b0b vdd b0a b3b b5a
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_1/dum0_in b0a b2b b1b b0b b0a b1b
+ b5b b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_1/out_5
+ b0b b2a rheo_3v_column_1/out_4 b4a b0b vdd b2b b0a b2b b0b vdd rheo_3v_column_1/res0_in
+ b0a b0a b1a b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_1/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_2 b5a b3a b0b b0b b2a rheo_3v_column_2/dum1_out b0b vdd b0a b3b b5b
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_2/dum0_in b0a b2b b1b b0b b0a b1b
+ b5a b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_3/out_5
+ b0b b2a rheo_3v_column_2/out_4 b4a b0b vdd b2b b0a b2b b0b vdd rheo_3v_column_2/res0_in
+ b0a b0a b1a b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_2/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_3 b5a b3a b0b b0b b2a rheo_3v_column_3/dum1_out b0b vdd b0a b3b b5a
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_3/dum0_in b0a b2b b1b b0b b0a b1b
+ b5b b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_3/out_5
+ b0b b2a rheo_3v_column_3/out_4 b4a b0b vdd b2b b0a b2b b0b vdd rheo_3v_column_3/res0_in
+ b0a b0a b1a b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_3/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_4 b5a b3a b0b b0b b2a rheo_3v_column_4/dum1_out b0b vdd b0a b3b b5b
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_4/dum0_in b0a b2b b1b b0b b0a b1b
+ b5a b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_5/out_5
+ b0b b2a rheo_3v_column_4/out_4 b4a b0b vdd b2b b0a b2b b0b vdd rheo_3v_column_4/res0_in
+ b0a b0a b1a b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_4/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_5 b5a b3a b0b b0b b2a rheo_3v_column_5/dum1_out b0b vdd b0a b3b b5a
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_5/dum0_in b0a b2b b1b b0b b0a b1b
+ b5b b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_5/out_5
+ b0b b2a rheo_3v_column_5/out_4 b4a b0b vdd b2b b0a b2b b0b vdd rheo_3v_column_5/res0_in
+ b0a b0a b1a b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_5/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_6 b5a b3a b0b b0b b2a rheo_3v_column_6/dum1_out b0b vdd b0a b3b b5b
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_6/dum0_in b0a b2b b1b b0b b0a b1b
+ b5a b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_7/out_5
+ b0b b2a rheo_3v_column_6/out_4 b4a b0b vdd b2b b0a b2b b0b vdd rheo_3v_column_6/res0_in
+ b0a b0a b1a b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_6/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_7 b5a b3a b0b b0b b2a rheo_3v_column_7/dum1_out b0b vdd b0a b3b b5a
+ b1b b0a vdd b0b b0a b1b vdd b0a rheo_3v_column_7/dum0_in b0a b2b b1b b0b b0a b1b
+ b5b b1b b1b b1b b3b b3a b1b b0a vdd b0b vdd vdd b0a b0a b0b b0a rheo_3v_column_7/out_5
+ b0b b2a rheo_3v_column_7/out_4 b4a b0b vdd b2b b0a b2b b0b vdd rheo_3v_column_7/res0_in
+ b0a b0a b1a b1a b1a b1a b4b b1a b2a b1a b1a vdd b2b b0a vdd b0b b0a b0b rheo_3v_column_7/res1_out
+ b0b b5b b0b b0a vdd b1a b0b b0b b2a vss rheo_3v_column
Xrheo_3v_column_odd_0 b5a b6b rheo_3v_column_0/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_2/in_5 b0a b3b b0a b0b b3a b1b b6a b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b rheo_3v_column_1/out_5 b1b
+ rheo_3v_column_0/dum1_out rheo_3v_column_1/res0_in vdd b2b b0a b1b b4b rheo_3v_column_0/out_4
+ b1a b2b b1b vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b
+ b1b vdd b0b rheo_3v_column_1/dum0_in b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b
+ b2a rheo_3v_column_odd
Xrheo_3v_column_odd_1 b5a b7b rheo_3v_column_1/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_2/in_5 b0a b3b b0a b0b b3a b1b b7a b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b out b1b rheo_3v_column_1/dum1_out
+ rheo_3v_column_2/res0_in vdd b2b b0a b1b b4b rheo_3v_column_1/out_4 b1a b2b b1b
+ vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b b1b vdd b0b
+ rheo_3v_column_2/dum0_in b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b b2a rheo_3v_column_odd
Xrheo_3v_column_odd_2 b5a b6a rheo_3v_column_2/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_2/in_5 b0a b3b b0a b0b b3a b1b b6b b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b rheo_3v_column_3/out_5 b1b
+ rheo_3v_column_2/dum1_out rheo_3v_column_3/res0_in vdd b2b b0a b1b b4b rheo_3v_column_2/out_4
+ b1a b2b b1b vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b
+ b1b vdd b0b rheo_3v_column_3/dum0_in b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b
+ b2a rheo_3v_column_odd
Xrheo_3v_column_odd_3 b5a vdd rheo_3v_column_3/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_3/in_5 b0a b3b b0a b0b b3a b1b vss b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b rheo_3v_column_odd_3/in_5
+ b1b rheo_3v_column_3/dum1_out rheo_3v_column_4/res0_in vdd b2b b0a b1b b4b rheo_3v_column_3/out_4
+ b1a b2b b1b vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b
+ b1b vdd b0b rheo_3v_column_4/dum0_in b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b
+ b2a rheo_3v_column_odd
Xrheo_3v_column_odd_4 b5a b6b rheo_3v_column_4/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_6/in_5 b0a b3b b0a b0b b3a b1b b6a b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b rheo_3v_column_5/out_5 b1b
+ rheo_3v_column_4/dum1_out rheo_3v_column_5/res0_in vdd b2b b0a b1b b4b rheo_3v_column_4/out_4
+ b1a b2b b1b vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b
+ b1b vdd b0b rheo_3v_column_5/dum0_in b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b
+ b2a rheo_3v_column_odd
Xrheo_3v_column_odd_5 b5a b7a rheo_3v_column_5/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_6/in_5 b0a b3b b0a b0b b3a b1b b7b b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b out b1b rheo_3v_column_5/dum1_out
+ rheo_3v_column_6/res0_in vdd b2b b0a b1b b4b rheo_3v_column_5/out_4 b1a b2b b1b
+ vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b b1b vdd b0b
+ rheo_3v_column_6/dum0_in b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b b2a rheo_3v_column_odd
Xrheo_3v_column_odd_6 b5a b6a rheo_3v_column_6/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_6/in_5 b0a b3b b0a b0b b3a b1b b6b b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b rheo_3v_column_7/out_5 b1b
+ rheo_3v_column_6/dum1_out rheo_3v_column_7/res0_in vdd b2b b0a b1b b4b rheo_3v_column_6/out_4
+ b1a b2b b1b vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b
+ b1b vdd b0b rheo_3v_column_7/dum0_in b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b
+ b2a rheo_3v_column_odd
Xrheo_3v_column_odd_7 b5a vdd rheo_3v_column_7/res1_out b0b b2a b0b b0b vdd b0a b1b
+ vdd b0b b0b b0a b1b rheo_3v_column_odd_7/in_5 b0a b3b b0a b0b b3a b1b vss b0b b0a
+ b2a b0b b0a vdd b0a vdd vdd b0a b0a b0a b3a b1b b4a b2b rheo_3v_column_odd_7/in_5
+ b1b rheo_3v_column_7/dum1_out Vlow vdd b2b b0a b1b b4b rheo_3v_column_7/out_4 b1a
+ b2b b1b vdd vdd vdd b1a b0a b0a b0b b2b b1a b1a b1a b0a b1a b1a b0b b2a b3b b1b
+ vdd b0b rheo_3v_column_odd_7/dum_out1 b0b b0a b0a b0b b5b b0b vdd b1a vss b0b b0b
+ b2a rheo_3v_column_odd
Xrheo_3v_column_dummy_0 b0a b1b b2a b1a b0b vss vdd b0a b0b vss vdd b0b b0a b0a b0b
+ b0a b0b b0b b0a vdd b0b b0a b2b b1a b0b b0a b0b vss vdd b0a vdd vdd vdd vss vdd
+ b0b vdd b0a b0b b4a b0a b0b b1a vdd b0a vdd b0b vdd b1b b0a vdd b2b vss vss b4b
+ vdd b1b b3a b1a b2b b2a b1a vdd b1a b1b vdd b3b b3a b1b b1a b2a b2b b1a b1b b3b
+ b5b vss vss b5a b1b b1b vdd vdd vdd b0a b0b Vhigh b0a b2a m1_6292_841# b0b rheo_3v_column_0/dum0_in
+ b0a b0b m1_6292_841# vss rheo_3v_column_dummy
Xrheo_3v_column_dummy_1 b0a b1b b2a b1a b0b vss vdd b0a b0b vss vdd b0b b0a b0a b0b
+ b0a b0b b0b b0a vdd b0b b0a b2b b1a b0b b0a b0b vss vdd b0a vdd vdd vdd vss vdd
+ b0b vdd b0a b0b b4a b0a b0b b1a vdd b0a vdd b0b vdd b1b b0a vdd b2b vss vss b4b
+ vdd b1b b3a b1a b2b b2a b1a vdd b1a b1b vdd b3b b3a b1b b1a b2a b2b b1a b1b b3b
+ b5b vss vss b5a b1b b1b vdd vdd vdd b0a b0b m1_25337_837# b0a b2a Vlow b0b m1_25337_837#
+ b0a b0b rheo_3v_column_odd_7/dum_out1 vss rheo_3v_column_dummy
Xrheo_level_shifter_array_0 b0 b3b b3a b4 b0a b4a b7a b1 b0b b5 b4b b7b b1b b5a b1a
+ b6 b2 b5b b6b b2b b2a b3 b7 dvdd vdd b6a dvss rheo_level_shifter_array
.ends

.subckt switch_array_14 dvdd left_hgbw_opamp_out right_instramp_out isolated_switch_xlarge_1[3|2]/off
+ analog1_connect[0] isolated_switch_xlarge_1[3|1]/on left_instramp_out right_hgbw_opamp_out
+ isolated_switch_xlarge_1[1|1]/on amuxbusA avdd dvss isolated_switch_xlarge_1[0|2]/on
+ isolated_switch_xlarge_1[3|0]/on isolated_switch_xlarge_1[2|1]/on isolated_switch_xlarge_1[1|0]/on
+ analog1 isolated_switch_xlarge_1[2|0]/on analog0 isolated_switch_xlarge_1[3|2]/on
+ analog1_core isolated_switch_xlarge_1[1|2]/on analog0_core isolated_switch_xlarge_1[1|2]/off
+ amuxbusB analog0_connect[0] isolated_switch_xlarge_1[2|2]/on analog0_connect[1]
+ isolated_switch_xlarge_1[0|1]/on isolated_switch_xlarge_1[3|1]/off isolated_switch_xlarge_1[2|2]/off
+ analog1_connect[1] isolated_switch_xlarge_1[1|1]/off isolated_switch_xlarge_1[0|0]/on
+ isolated_switch_xlarge_1[0|2]/off isolated_switch_xlarge_1[3|0]/off isolated_switch_xlarge_1[2|0]/off
+ isolated_switch_xlarge_1[2|1]/off isolated_switch_xlarge_1[1|0]/off isolated_switch_xlarge_1[0|1]/off
+ right_lp_opamp_out isolated_switch_xlarge_1[0|0]/off left_lp_opamp_out avss
Xisolated_switch_xlarge_0[0] analog1_connect[0] analog1 analog1_core avdd analog1_connect[1]
+ avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_0[1] analog0_connect[0] analog0 analog0_core avdd analog0_connect[1]
+ avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_1[0|0] isolated_switch_xlarge_1[0|0]/on right_lp_opamp_out
+ amuxbusB avdd isolated_switch_xlarge_1[0|0]/off avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_1[1|0] isolated_switch_xlarge_1[1|0]/on right_lp_opamp_out
+ analog1_core avdd isolated_switch_xlarge_1[1|0]/off avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_1[2|0] isolated_switch_xlarge_1[2|0]/on right_instramp_out
+ amuxbusA avdd isolated_switch_xlarge_1[2|0]/off avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_1[3|0] isolated_switch_xlarge_1[3|0]/on right_instramp_out
+ analog0_core avdd isolated_switch_xlarge_1[3|0]/off avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_1[0|1] isolated_switch_xlarge_1[0|1]/on left_hgbw_opamp_out
+ amuxbusB avdd isolated_switch_xlarge_1[0|1]/off avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_1[1|1] isolated_switch_xlarge_1[1|1]/on left_hgbw_opamp_out
+ analog1_core avdd isolated_switch_xlarge_1[1|1]/off avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_1[2|1] isolated_switch_xlarge_1[2|1]/on right_hgbw_opamp_out
+ amuxbusA avdd isolated_switch_xlarge_1[2|1]/off avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_1[3|1] isolated_switch_xlarge_1[3|1]/on right_hgbw_opamp_out
+ analog0_core avdd isolated_switch_xlarge_1[3|1]/off avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_1[0|2] isolated_switch_xlarge_1[0|2]/on left_instramp_out
+ amuxbusB avdd isolated_switch_xlarge_1[0|2]/off avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_1[1|2] isolated_switch_xlarge_1[1|2]/on left_instramp_out
+ analog1_core avdd isolated_switch_xlarge_1[1|2]/off avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_1[2|2] isolated_switch_xlarge_1[2|2]/on left_lp_opamp_out
+ amuxbusA avdd isolated_switch_xlarge_1[2|2]/off avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_1[3|2] isolated_switch_xlarge_1[3|2]/on left_lp_opamp_out
+ analog0_core avdd isolated_switch_xlarge_1[3|2]/off avss dvdd dvss isolated_switch_xlarge
.ends

.subckt simple_switch_array_6 simplest_analog_switch_ena1v8_1[0]/in simplest_analog_switch_ena1v8_0[2]/in
+ simplest_analog_switch_ena1v8_0[0]/in simplest_analog_switch_ena1v8_0[2]/out simplest_analog_switch_ena1v8_1[2]/on
+ simplest_analog_switch_ena1v8_1[1]/on simplest_analog_switch_ena1v8_1[0]/on simplest_analog_switch_ena1v8_0[2]/on
+ simplest_analog_switch_ena1v8_1[2]/in simplest_analog_switch_ena1v8_1[2]/avdd simplest_analog_switch_ena1v8_1[1]/in
+ simplest_analog_switch_ena1v8_1[2]/dvdd simplest_analog_switch_ena1v8_1[2]/out simplest_analog_switch_ena1v8_0[0]/on
+ simplest_analog_switch_ena1v8_0[1]/in simplest_analog_switch_ena1v8_0[1]/on simplest_analog_switch_ena1v8_1[2]/avss
+ VSUBS
Xsimplest_analog_switch_ena1v8_0[0] simplest_analog_switch_ena1v8_1[2]/avdd simplest_analog_switch_ena1v8_1[2]/dvdd
+ simplest_analog_switch_ena1v8_1[2]/avss simplest_analog_switch_ena1v8_0[0]/on simplest_analog_switch_ena1v8_0[2]/out
+ VSUBS simplest_analog_switch_ena1v8_0[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[1] simplest_analog_switch_ena1v8_1[2]/avdd simplest_analog_switch_ena1v8_1[2]/dvdd
+ simplest_analog_switch_ena1v8_1[2]/avss simplest_analog_switch_ena1v8_0[1]/on simplest_analog_switch_ena1v8_0[2]/out
+ VSUBS simplest_analog_switch_ena1v8_0[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[2] simplest_analog_switch_ena1v8_1[2]/avdd simplest_analog_switch_ena1v8_1[2]/dvdd
+ simplest_analog_switch_ena1v8_1[2]/avss simplest_analog_switch_ena1v8_0[2]/on simplest_analog_switch_ena1v8_0[2]/out
+ VSUBS simplest_analog_switch_ena1v8_0[2]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[0] simplest_analog_switch_ena1v8_1[2]/avdd simplest_analog_switch_ena1v8_1[2]/dvdd
+ simplest_analog_switch_ena1v8_1[2]/avss simplest_analog_switch_ena1v8_1[0]/on simplest_analog_switch_ena1v8_1[2]/out
+ VSUBS simplest_analog_switch_ena1v8_1[0]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1] simplest_analog_switch_ena1v8_1[2]/avdd simplest_analog_switch_ena1v8_1[2]/dvdd
+ simplest_analog_switch_ena1v8_1[2]/avss simplest_analog_switch_ena1v8_1[1]/on simplest_analog_switch_ena1v8_1[2]/out
+ VSUBS simplest_analog_switch_ena1v8_1[1]/in simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[2] simplest_analog_switch_ena1v8_1[2]/avdd simplest_analog_switch_ena1v8_1[2]/dvdd
+ simplest_analog_switch_ena1v8_1[2]/avss simplest_analog_switch_ena1v8_1[2]/on simplest_analog_switch_ena1v8_1[2]/out
+ VSUBS simplest_analog_switch_ena1v8_1[2]/in simplest_analog_switch_ena1v8
.ends

.subckt sky130_fd_pr__nfet_01v8_QXBCRM a_n1000_n188# a_n1160_n274# a_1000_n100# a_n1058_n100#
X0 a_1000_n100# a_n1000_n188# a_n1058_n100# a_n1160_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_B5H3CA w_n1196_n319# a_n1000_n197# a_1000_n100#
+ a_n1058_n100#
X0 a_1000_n100# a_n1000_n197# a_n1058_n100# w_n1196_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
.ends

.subckt buffer input output vbias vss vdd
XXM1 input vss m1_2942_n986# m1_772_n974# sky130_fd_pr__nfet_01v8_QXBCRM
XXM2 output vss output m1_2942_n986# sky130_fd_pr__nfet_01v8_QXBCRM
XXM3 vdd m1_772_n974# vdd m1_772_n974# sky130_fd_pr__pfet_01v8_lvt_B5H3CA
XXM4 vdd m1_772_n974# output vdd sky130_fd_pr__pfet_01v8_lvt_B5H3CA
XXM5 vbias vss m1_2942_n986# vss sky130_fd_pr__nfet_01v8_QXBCRM
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__0 a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base m=1
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_3VR9VM w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_6VRZAW a_100_n536# w_n296_n1191# a_n100_675# a_100_336#
+ a_n158_n536# a_n158_772# a_n100_n633# a_n100_239# a_n100_n197# a_100_n100# a_n158_336#
+ a_100_n972# a_n158_n100# a_100_772# a_n158_n972# a_n100_n1069#
X0 a_100_336# a_n100_239# a_n158_336# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 a_100_772# a_n100_675# a_n158_772# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_100_n536# a_n100_n633# a_n158_n536# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X4 a_100_n972# a_n100_n1069# a_n158_n972# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_3HMWVM w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_69TQ3K a_n260_n274# a_100_n100# a_n158_n100# a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n260_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_od_ip__tempsensor_ext_vp vbe2_out vbe1_out ena vbg vdd vss
Xx1 x1/input vbe2_out ena vss vdd buffer
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RJ_1 vss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__0
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0 vss vbg sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__0
Xx2 x2/input vbe1_out ena vss vdd buffer
XXQ_BR1 x1/input vss vss sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
XXQ_BL1 x2/input vss vss sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
XXM11 vdd vp vdd x2/input sky130_fd_pr__pfet_01v8_lvt_3VR9VM
XXM22 vdd vdd vp vdd x1/input x1/input vp vp vp vdd x1/input vdd x1/input vdd x1/input
+ vp sky130_fd_pr__pfet_01v8_lvt_6VRZAW
XXM33 vdd ena vp vdd sky130_fd_pr__pfet_01v8_3HMWVM
XXM44 vss m1_772_n1144# m1_420_n380# vbg sky130_fd_pr__nfet_01v8_69TQ3K
XXM55 vss vp m1_772_n1144# vp sky130_fd_pr__nfet_01v8_69TQ3K
XXM66 ena vss m1_772_n1144# vss sky130_fd_pr__nfet_01v8_QXBCRM
XXM77 vdd m1_420_n380# vp vdd sky130_fd_pr__pfet_01v8_3HMWVM
XXM88 vdd m1_420_n380# vdd m1_420_n380# sky130_fd_pr__pfet_01v8_3HMWVM
.ends

.subckt switch_array_2 channel0_in_to_out[1] channel0_in_to_out[0] channel1_in_to_out[1]
+ channel1_in_to_out[0] channel0_in channel1_in channel1_out avdd dvss channel0_out
+ dvdd avss
Xisolated_switch_xlarge_0[0] channel1_in_to_out[0] channel1_out channel1_in avdd channel1_in_to_out[1]
+ avss dvdd dvss isolated_switch_xlarge
Xisolated_switch_xlarge_0[1] channel0_in_to_out[0] channel0_out channel0_in avdd channel0_in_to_out[1]
+ avss dvdd dvss isolated_switch_xlarge
.ends

.subckt simple_analog_mux_sel1v8 inA out avdd dvdd selA inB dvss avss
Xsimple_analog_switch_2_0 sky130_fd_sc_hvl__inv_2_0/Y avdd avss sky130_fd_sc_hvl__inv_2_1/Y
+ out inA simple_analog_switch_2
Xsimple_analog_switch_2_1 sky130_fd_sc_hvl__inv_2_1/Y avdd avss sky130_fd_sc_hvl__inv_2_0/Y
+ inB out simple_analog_switch_2
Xsky130_fd_sc_hvl__inv_2_0 sky130_fd_sc_hvl__inv_2_1/Y dvss dvss avdd avdd sky130_fd_sc_hvl__inv_2_0/Y
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_1 sky130_fd_sc_hvl__inv_2_1/A dvss dvss avdd avdd sky130_fd_sc_hvl__inv_2_1/Y
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 selA dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_1/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__diode_2_0 selA dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_0 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__decap_4_1 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_4V4BDM a_n29_n50# a_n187_n50# w_n387_n347# a_29_n147#
+ a_n129_n147# a_129_n50#
X0 a_129_n50# a_29_n147# a_n29_n50# w_n387_n347# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1 a_n29_n50# a_n129_n147# a_n187_n50# w_n387_n347# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_8T5BGA a_n187_n136# a_129_n136# w_n387_n362#
+ a_29_n162# a_n129_n162# a_n29_n136#
X0 a_n29_n136# a_n129_n162# a_n187_n136# w_n387_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X1 a_129_n136# a_29_n162# a_n29_n136# w_n387_n362# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_C5EREZ a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_S48KL6 a_n321_n322# a_n29_n100# a_n187_n100#
+ a_129_n100# a_29_n188# a_n129_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n188# a_n187_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt level_shifter_up VDD_HV x_lv x_hv xb_hv VDD_LV VSUBS m1_380_440# GND_HV
Xsky130_fd_pr__pfet_g5v0d10v5_4V4BDM_0 VDD_HV xb_hv VDD_HV xb_hv x_hv x_hv sky130_fd_pr__pfet_g5v0d10v5_4V4BDM
Xsky130_fd_pr__pfet_g5v0d10v5_8T5BGA_0 m1_380_440# m1_380_440# VDD_LV x_lv x_lv VDD_LV
+ sky130_fd_pr__pfet_g5v0d10v5_8T5BGA
Xsky130_fd_pr__nfet_g5v0d10v5_C5EREZ_0 m1_380_440# VSUBS VSUBS x_lv sky130_fd_pr__nfet_g5v0d10v5_C5EREZ
Xsky130_fd_pr__nfet_g5v0d10v5_S48KL6_0 GND_HV GND_HV x_hv xb_hv x_lv m1_380_440# sky130_fd_pr__nfet_g5v0d10v5_S48KL6
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_RUG6CB a_n400_n497# a_400_n400# w_n658_n697#
+ a_n458_n400#
X0 a_400_n400# a_n400_n497# a_n458_n400# w_n658_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=4
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_M7X63G a_150_n800# a_n208_n800# a_n150_n888#
+ a_n342_n1022#
X0 a_150_n800# a_n150_n888# a_n208_n800# a_n342_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_REE66T a_n487_n497# a_487_n400# a_n29_n400# a_545_n497#
+ a_n803_n400# a_29_n497# a_n287_n400# a_n1061_n400# a_n745_n497# a_803_n497# a_745_n400#
+ a_n229_n497# a_287_n497# a_n1003_n497# a_229_n400# a_n545_n400# w_n1261_n697# a_1003_n400#
X0 a_n545_n400# a_n745_n497# a_n803_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X1 a_n803_n400# a_n1003_n497# a_n1061_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X2 a_n287_n400# a_n487_n497# a_n545_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 a_1003_n400# a_803_n497# a_745_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X4 a_487_n400# a_287_n497# a_229_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X5 a_745_n400# a_545_n497# a_487_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X6 a_229_n400# a_29_n497# a_n29_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X7 a_n29_n400# a_n229_n497# a_n287_n400# w_n1261_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_LUSSBJ a_108_n288# a_50_n200# a_n208_n288# a_n400_n422#
+ a_n108_n200# a_n266_n200# a_n50_n288# a_208_n200#
X0 a_n108_n200# a_n208_n288# a_n266_n200# a_n400_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X1 a_208_n200# a_108_n288# a_50_n200# a_n400_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2 a_50_n200# a_n50_n288# a_n108_n200# a_n400_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__res_high_po_2p85_EP2UD7 a_n2283_n3624# a_381_n3624# a_n2437_n3778#
+ a_n285_3192# a_1047_3192# a_n951_3192# a_1713_3192# a_n1617_n3624# a_381_3192# a_n285_n3624#
+ a_n951_n3624# a_1047_n3624# a_n2283_3192# a_1713_n3624# a_n1617_3192#
X0 a_n285_3192# a_n285_n3624# a_n2437_n3778# sky130_fd_pr__res_high_po_2p85 l=32.08
X1 a_1047_3192# a_1047_n3624# a_n2437_n3778# sky130_fd_pr__res_high_po_2p85 l=32.08
X2 a_n951_3192# a_n951_n3624# a_n2437_n3778# sky130_fd_pr__res_high_po_2p85 l=32.08
X3 a_1713_3192# a_1713_n3624# a_n2437_n3778# sky130_fd_pr__res_high_po_2p85 l=32.08
X4 a_n2283_3192# a_n2283_n3624# a_n2437_n3778# sky130_fd_pr__res_high_po_2p85 l=32.08
X5 a_n1617_3192# a_n1617_n3624# a_n2437_n3778# sky130_fd_pr__res_high_po_2p85 l=32.08
X6 a_381_3192# a_381_n3624# a_n2437_n3778# sky130_fd_pr__res_high_po_2p85 l=32.08
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TAUUP3 a_n345_n431# a_129_n431# a_29_n457# a_n129_n457#
+ a_287_n431# a_187_n457# a_n287_n457# a_n29_n431# a_n479_n591# a_n187_n431#
X0 a_n187_n431# a_n287_n457# a_n345_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_287_n431# a_187_n457# a_129_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2 a_129_n431# a_29_n457# a_n29_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n29_n431# a_n129_n457# a_n187_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_RJSTGP a_29_n297# a_n887_n200# a_n29_n200# a_n829_n297#
+ w_n1087_n497# a_829_n200#
X0 a_n29_n200# a_n829_n297# a_n887_n200# w_n1087_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=4
X1 a_829_n200# a_29_n297# a_n29_n200# w_n1087_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=4
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_8JQF8T a_n100_n1015# a_n158_118# a_n100_21# w_n358_n1215#
+ a_100_n918# a_n158_n918# a_100_118#
X0 a_100_118# a_n100_21# a_n158_118# w_n358_n1215# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X1 a_100_n918# a_n100_n1015# a_n158_n918# w_n358_n1215# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_MMHSE7 a_100_n400# a_n292_n622# a_n158_n400#
+ a_n100_n488#
X0 a_100_n400# a_n100_n488# a_n158_n400# a_n292_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_PNRDLC a_n150_n897# a_150_n800# w_n408_n1097#
+ a_n208_n800#
X0 a_150_n800# a_n150_n897# a_n208_n800# w_n408_n1097# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_46Z5PG a_129_n200# a_29_n288# a_n129_n288# a_n321_n422#
+ a_n29_n200# a_n187_n200#
X0 a_129_n200# a_29_n288# a_n29_n200# a_n321_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X1 a_n29_n200# a_n129_n288# a_n187_n200# a_n321_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_RRA4TL a_n258_n50# a_n200_n138# a_200_n50# a_n392_n272#
X0 a_200_n50# a_n200_n138# a_n258_n50# a_n392_n272# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CRL9SD a_n150_n897# a_150_n800# w_n408_n1097#
+ a_n208_n800#
X0 a_150_n800# a_n150_n897# a_n208_n800# w_n408_n1097# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1.5
.ends

.subckt sky130_fd_pr__pfet_01v8_YTEHH6 w_n425_n619# a_n29_n400# a_29_n497# a_n287_n400#
+ a_n229_n497# a_229_n400#
X0 a_n29_n400# a_n229_n497# a_n287_n400# w_n425_n619# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X1 a_229_n400# a_29_n497# a_n29_n400# w_n425_n619# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_8TUSME a_n345_n200# a_129_n200# a_287_n200# a_n479_n422#
+ a_29_n288# a_n129_n288# a_187_n288# a_n287_n288# a_n29_n200# a_n187_n200#
X0 a_n187_n200# a_n287_n288# a_n345_n200# a_n479_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X1 a_287_n200# a_187_n288# a_129_n200# a_n479_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2 a_129_n200# a_29_n288# a_n29_n200# a_n479_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X3 a_n29_n200# a_n129_n288# a_n187_n200# a_n479_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_T8W2FW a_150_n800# a_n208_n800# a_n150_n888#
+ a_n342_n1022#
X0 a_150_n800# a_n150_n888# a_n208_n800# a_n342_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_AUB4P8 a_150_n800# a_n208_n800# a_n150_n888#
+ a_n342_n1022#
X0 a_150_n800# a_n150_n888# a_n208_n800# a_n342_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1.5
.ends

.subckt sky130_fd_pr__nfet_01v8_HWT53N a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_LHNF5N a_n345_n431# a_129_n431# a_29_n457# a_n129_n457#
+ a_287_n431# a_187_n457# a_n287_n457# a_n29_n431# a_n479_n591# a_n187_n431#
X0 a_n187_n431# a_n287_n457# a_n345_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_287_n431# a_187_n457# a_129_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2 a_129_n431# a_29_n457# a_n29_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n29_n431# a_n129_n457# a_n187_n431# a_n479_n591# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_EPRAC4 a_15_n200# w_n211_n419# a_n33_n297# a_n73_n200#
X0 a_15_n200# a_n33_n297# a_n73_n200# w_n211_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Q8UPKT a_n829_n615# w_n1087_n815# a_29_n615#
+ a_29_21# a_n887_n518# a_829_118# a_n29_n518# a_829_n518# a_n29_118# a_n887_118#
+ a_n829_21#
X0 a_829_118# a_29_21# a_n29_118# w_n1087_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=4
X1 a_n29_118# a_n829_21# a_n887_118# w_n1087_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=4
X2 a_n29_n518# a_n829_n615# a_n887_n518# w_n1087_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=4
X3 a_829_n518# a_29_n615# a_n29_n518# w_n1087_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=4
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_MRHAE7 a_100_n400# a_n292_n622# a_n158_n400#
+ a_n100_n488#
X0 a_100_n400# a_n100_n488# a_n158_n400# a_n292_n622# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_X332GA a_29_n297# a_n129_n297# a_129_n200# a_n29_n200#
+ w_n387_n497# a_n187_n200#
X0 a_129_n200# a_29_n297# a_n29_n200# w_n387_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X1 a_n29_n200# a_n129_n297# a_n187_n200# w_n387_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_4RA4DJ a_n603_n288# a_n345_n200# a_129_n200#
+ a_n503_n200# a_287_n200# a_n661_n200# a_445_n200# a_29_n288# a_n129_n288# a_603_n200#
+ a_187_n288# a_n795_n422# a_n287_n288# a_345_n288# a_n29_n200# a_n187_n200# a_n445_n288#
+ a_503_n288#
X0 a_n187_n200# a_n287_n288# a_n345_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X1 a_287_n200# a_187_n288# a_129_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X2 a_n345_n200# a_n445_n288# a_n503_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X3 a_129_n200# a_29_n288# a_n29_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X4 a_445_n200# a_345_n288# a_287_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X5 a_n503_n200# a_n603_n288# a_n661_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X6 a_n29_n200# a_n129_n288# a_n187_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X7 a_603_n200# a_503_n288# a_445_n200# a_n795_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_GHE6BF a_n158_n518# a_n158_118# a_n100_21# a_n100_n615#
+ w_n358_n815# a_100_118# a_100_n518#
X0 a_100_118# a_n100_21# a_n158_118# w_n358_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X1 a_100_n518# a_n100_n615# a_n158_n518# w_n358_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WGHV7X a_400_n509# a_n458_109# a_n400_21# a_n458_n509#
+ a_n592_n731# a_400_109# a_n400_n597#
X0 a_400_n509# a_n400_n597# a_n458_n509# a_n592_n731# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
X1 a_400_109# a_n400_21# a_n458_109# a_n592_n731# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_LURNA9 a_n287_n200# a_n1061_n200# a_745_n200#
+ a_n487_n288# a_545_n288# a_229_n200# a_n1195_n422# a_n545_n200# a_29_n288# a_n745_n288#
+ a_1003_n200# a_803_n288# a_487_n200# a_n29_n200# a_n229_n288# a_287_n288# a_n1003_n288#
+ a_n803_n200#
X0 a_n29_n200# a_n229_n288# a_n287_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_229_n200# a_29_n288# a_n29_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_n545_n200# a_n745_n288# a_n803_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_n803_n200# a_n1003_n288# a_n1061_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X4 a_n287_n200# a_n487_n288# a_n545_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_745_n200# a_545_n288# a_487_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_1003_n200# a_803_n288# a_745_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X7 a_487_n200# a_287_n288# a_229_n200# a_n1195_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_RM8L2M a_n258_n50# a_n200_n138# a_200_n50# a_n392_n272#
X0 a_200_n50# a_n200_n138# a_n258_n50# a_n392_n272# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_N8ANR9 a_n345_n364# a_129_n364# a_287_n364# w_n545_n662#
+ a_29_n461# a_n129_n461# a_187_n461# a_n287_n461# a_n29_n364# a_n187_n364#
X0 a_n187_n364# a_n287_n461# a_n345_n364# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 a_287_n364# a_187_n461# a_129_n364# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2 a_129_n364# a_29_n461# a_n29_n364# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n29_n364# a_n129_n461# a_n187_n364# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CDNABP a_n100_n597# a_n100_21# a_100_109# a_100_n509#
+ a_n158_n509# a_n292_n731# a_n158_109#
X0 a_100_n509# a_n100_n597# a_n158_n509# a_n292_n731# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X1 a_100_109# a_n100_21# a_n158_109# a_n292_n731# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_6UJQA2 a_n187_n436# a_n345_n436# a_129_n436#
+ a_287_n436# w_n545_n662# a_29_n462# a_n129_n462# a_187_n462# a_n287_n462# a_n29_n436#
X0 a_129_n436# a_29_n462# a_n29_n436# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X1 a_n29_n436# a_n129_n462# a_n187_n436# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 a_n187_n436# a_n287_n462# a_n345_n436# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X3 a_287_n436# a_187_n462# a_129_n436# w_n545_n662# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CS979Q a_n400_n615# a_400_118# w_n658_n815# a_n400_21#
+ a_400_n518# a_n458_118# a_n458_n518#
X0 a_400_118# a_n400_21# a_n458_118# w_n658_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
X1 a_400_n518# a_n400_n615# a_n458_n518# w_n658_n815# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_2CKAKF a_n819_n200# a_n345_n200# a_n977_n200#
+ a_n1135_n200# a_29_n297# a_n129_n297# a_187_n297# a_129_n200# a_n503_n200# a_n1293_n200#
+ a_n287_n297# a_819_n297# a_345_n297# a_n1077_n297# a_287_n200# a_n661_n200# a_n919_n297#
+ a_977_n297# a_n445_n297# a_919_n200# a_503_n297# a_n1235_n297# a_445_n200# a_1135_n297#
+ a_n603_n297# a_1077_n200# a_661_n297# a_603_n200# w_n1493_n497# a_n761_n297# a_1235_n200#
+ a_761_n200# a_n29_n200# a_n187_n200#
X0 a_n819_n200# a_n919_n297# a_n977_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X1 a_n661_n200# a_n761_n297# a_n819_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X2 a_919_n200# a_819_n297# a_761_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X3 a_n187_n200# a_n287_n297# a_n345_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X4 a_761_n200# a_661_n297# a_603_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X5 a_287_n200# a_187_n297# a_129_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X6 a_n345_n200# a_n445_n297# a_n503_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X7 a_129_n200# a_29_n297# a_n29_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X8 a_445_n200# a_345_n297# a_287_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X9 a_n977_n200# a_n1077_n297# a_n1135_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X10 a_n503_n200# a_n603_n297# a_n661_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X11 a_1077_n200# a_977_n297# a_919_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X12 a_n29_n200# a_n129_n297# a_n187_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X13 a_603_n200# a_503_n297# a_445_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X14 a_1235_n200# a_1135_n297# a_1077_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X15 a_n1135_n200# a_n1235_n297# a_n1293_n200# w_n1493_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EEFBWQ a_400_n200# a_n592_n422# a_n458_n200#
+ a_n400_n288#
X0 a_400_n200# a_n400_n288# a_n458_n200# a_n592_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_9432CF a_n345_n200# a_29_n297# a_n129_n297# w_n703_n497#
+ a_187_n297# a_129_n200# a_n503_n200# a_n287_n297# a_345_n297# a_287_n200# a_n445_n297#
+ a_445_n200# a_n29_n200# a_n187_n200#
X0 a_n187_n200# a_n287_n297# a_n345_n200# w_n703_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X1 a_287_n200# a_187_n297# a_129_n200# w_n703_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X2 a_n345_n200# a_n445_n297# a_n503_n200# w_n703_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X3 a_129_n200# a_29_n297# a_n29_n200# w_n703_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X4 a_445_n200# a_345_n297# a_287_n200# w_n703_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X5 a_n29_n200# a_n129_n297# a_n187_n200# w_n703_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_2432J2 a_n345_n200# a_29_n297# a_n129_n297# a_187_n297#
+ a_129_n200# a_n287_n297# a_287_n200# a_n29_n200# a_n187_n200# w_n545_n497#
X0 a_n187_n200# a_n287_n297# a_n345_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X1 a_287_n200# a_187_n297# a_129_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2 a_129_n200# a_29_n297# a_n29_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X3 a_n29_n200# a_n129_n297# a_n187_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_ak_ip__comparator Vinp Vinm AVDD en hyst[1] hyst[0] trim[5] trim[4]
+ trim[3] trim[2] trim[1] trim[0] Vout DVDD ibias DGND AGND
Xlevel_shifter_up_3 AVDD en en_hv enb_hv DVDD DGND m1_36128_n32592# AGND level_shifter_up
Xsky130_fd_pr__pfet_g5v0d10v5_RUG6CB_0 m1_25710_11400# AVDD AVDD m1_25710_11400# sky130_fd_pr__pfet_g5v0d10v5_RUG6CB
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_60 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_82 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_REE66T_1 m1_36250_n26840# m1_2500_n30560# m1_2500_n30560#
+ m1_36250_n26840# m1_31820_n13600# m1_36250_n26840# m1_31820_n13600# m1_2500_n30560#
+ m1_36250_n26840# m1_36250_n26840# m1_31820_n13600# m1_36250_n26840# m1_36250_n26840#
+ m1_36250_n26840# m1_31820_n13600# m1_2500_n30560# AVDD m1_2500_n30560# sky130_fd_pr__pfet_g5v0d10v5_REE66T
Xlevel_shifter_up_4 AVDD trim[3] level_shifter_up_4/x_hv trim3b_hv DVDD DGND m1_35128_n32592#
+ AGND level_shifter_up
Xsky130_fd_pr__nfet_g5v0d10v5_LUSSBJ_0 hyst0_hv AGND hyst0_hv AGND m1_33660_n1540#
+ AGND hyst0_hv m1_33660_n1540# sky130_fd_pr__nfet_g5v0d10v5_LUSSBJ
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_50 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_61 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_83 m1_420_6500# m1_2500_5340# m1_4100_9160# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__res_high_po_2p85_EP2UD7_0 AGND m1_25040_4590# AGND m1_24380_11400#
+ m1_25710_11400# m1_23050_11400# AGND m1_23040_4590# m1_24380_11400# m1_23710_4590#
+ m1_23710_4590# m1_25040_4590# AGND AGND m1_23050_11400# sky130_fd_pr__res_high_po_2p85_EP2UD7
Xlevel_shifter_up_5 AVDD trim[4] level_shifter_up_5/x_hv trim4b_hv DVDD DGND m1_34128_n32592#
+ AGND level_shifter_up
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_40 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_51 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_62 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_73 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_84 m1_420_6500# m1_2500_6140# m1_4100_8360# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__res_high_po_2p85_EP2UD7_1 AGND m1_24360_n31900# AGND m1_23690_n25080#
+ m1_25020_n25080# m1_23690_n25080# AGND m1_23030_n31900# m1_25020_n25080# m1_24360_n31900#
+ m1_23030_n31900# res_p_bot AGND AGND m1_23030_n25080# sky130_fd_pr__res_high_po_2p85_EP2UD7
Xlevel_shifter_up_6 AVDD trim[0] level_shifter_up_6/x_hv level_shifter_up_6/xb_hv
+ DVDD DGND level_shifter_up_6/m1_380_440# AGND level_shifter_up
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_30 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_41 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_52 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_63 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_74 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_85 m1_420_6500# m1_2500_6140# m1_4100_8360# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xlevel_shifter_up_7 AVDD trim[2] level_shifter_up_7/x_hv level_shifter_up_7/xb_hv
+ DVDD DGND level_shifter_up_7/m1_380_440# AGND level_shifter_up
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_20 m1_420_6500# m1_2500_6140# m1_4100_8360# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_31 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_42 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_53 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_75 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_86 m1_420_6500# m1_2500_5340# m1_4100_9160# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xlevel_shifter_up_8 AVDD trim[1] level_shifter_up_8/x_hv level_shifter_up_8/xb_hv
+ DVDD DGND level_shifter_up_8/m1_380_440# AGND level_shifter_up
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_10 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_21 m1_420_6500# m1_2500_6140# m1_4100_8360# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_32 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_43 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_54 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_76 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_87 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_11 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_22 m1_420_6500# m1_2500_5340# m1_4100_9160# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_33 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_44 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_55 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_77 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_88 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_12 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_23 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_34 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_45 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_78 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_TAUUP3_0 bias_n AGND enb_hv enb_hv bias_n enb_hv enb_hv
+ bias_n AGND AGND sky130_fd_pr__nfet_g5v0d10v5_TAUUP3
Xsky130_fd_pr__pfet_g5v0d10v5_RJSTGP_0 m1_29940_7140# AVDD m1_29940_7140# m1_29940_7140#
+ AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_RJSTGP
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_13 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_35 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_46 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_57 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_79 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_8JQF8T_0 Vop m1_29860_5120# Vom AVDD m1_29880_4800#
+ m1_29860_5120# m1_30900_4740# sky130_fd_pr__pfet_g5v0d10v5_8JQF8T
Xsky130_fd_pr__nfet_g5v0d10v5_MMHSE7_0 m1_29880_4800# AGND AGND m1_29880_4800# sky130_fd_pr__nfet_g5v0d10v5_MMHSE7
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_14 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_25 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_36 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_58 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_30 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_MMHSE7_1 DGND DGND m1_35390_11200# m1_29880_4800# sky130_fd_pr__nfet_g5v0d10v5_MMHSE7
Xsky130_fd_pr__nfet_g5v0d10v5_46Z5PG_0 AGND level_shifter_up_8/x_hv level_shifter_up_8/x_hv
+ AGND m1_32060_2060# AGND sky130_fd_pr__nfet_g5v0d10v5_46Z5PG
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_15 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_26 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_37 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_59 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_31 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_20 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_RRA4TL_0 m1_29880_4800# m1_30900_4740# AGND AGND sky130_fd_pr__nfet_g5v0d10v5_RRA4TL
Xsky130_fd_pr__nfet_g5v0d10v5_46Z5PG_1 AGND level_shifter_up_6/x_hv level_shifter_up_6/x_hv
+ AGND m1_35270_2060# AGND sky130_fd_pr__nfet_g5v0d10v5_46Z5PG
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_27 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_38 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_49 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_32 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_21 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_10 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|0] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|0] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|0] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|0] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|0] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|0] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|0] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|0] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|1] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|1] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|1] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|1] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|1] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|1] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|1] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|1] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|2] m1_4100_n29230# Vfold_bot_m AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|2] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|2] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|2] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|2] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|2] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|2] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|2] m1_4100_n29230# Vfold_bot_m AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|3] m1_4100_n28430# m1_2500_n30560# AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|3] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|3] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|3] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|3] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|3] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|3] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|3] m1_4100_n28430# m1_2500_n30560# AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|4] m1_4100_n28430# m1_2500_n30560# AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|4] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|4] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|4] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|4] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|4] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|4] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|4] m1_4100_n28430# m1_2500_n30560# AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|5] m1_4100_n29230# Vfold_bot_m AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|5] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|5] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|5] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|5] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|5] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|5] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|5] m1_4100_n29230# Vfold_bot_m AVDD m1_420_n29120#
+ sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|6] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|6] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|6] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|6] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|6] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|6] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|6] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|6] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[0|7] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[1|7] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[2|7] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[3|7] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[4|7] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[5|7] Vinm m1_2500_n30560# AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[6|7] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_g5v0d10v5_CRL9SD_0[7|7] Vinp Vfold_bot_m AVDD Vxp sky130_fd_pr__pfet_g5v0d10v5_CRL9SD
Xsky130_fd_pr__pfet_01v8_YTEHH6_0 DVDD m1_35390_11200# m1_35390_11200# DVDD m1_35390_11200#
+ DVDD sky130_fd_pr__pfet_01v8_YTEHH6
Xsky130_fd_pr__nfet_g5v0d10v5_8TUSME_0 DGND m1_35900_10510# DGND DGND enb_hv enb_hv
+ enb_hv enb_hv DGND m1_35900_10510# sky130_fd_pr__nfet_g5v0d10v5_8TUSME
Xsky130_fd_pr__nfet_g5v0d10v5_46Z5PG_2 AGND level_shifter_up_8/x_hv level_shifter_up_8/x_hv
+ AGND m1_32060_2060# AGND sky130_fd_pr__nfet_g5v0d10v5_46Z5PG
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_17 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_28 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_33 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_22 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_11 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_01v8_YTEHH6_1 DVDD m1_35900_10510# m1_35390_11200# DVDD m1_35390_11200#
+ DVDD sky130_fd_pr__pfet_01v8_YTEHH6
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_30 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_AUB4P8_0 m1_9080_4100# m1_7790_4530# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_AUB4P8
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_18 Vxm m1_2500_6140# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_29 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_34 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_23 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_12 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_31 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_20 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_01v8_HWT53N_0 DGND m1_35900_10510# m1_34800_n26840# DGND sky130_fd_pr__nfet_01v8_HWT53N
Xsky130_fd_pr__nfet_g5v0d10v5_AUB4P8_1 m1_9080_4100# m1_7790_4530# Vinm AGND sky130_fd_pr__nfet_g5v0d10v5_AUB4P8
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_19 m1_420_6500# m1_2500_5340# m1_4100_9160# AGND
+ sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_35 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_24 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_13 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_32 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_21 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_10 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_01v8_HWT53N_1 DGND m1_36250_n26840# Vout DGND sky130_fd_pr__nfet_01v8_HWT53N
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_9 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__nfet_g5v0d10v5_LHNF5N_0 m1_23030_n25080# m1_4100_n29230# trim5b_hv
+ trim5b_hv m1_23030_n25080# trim5b_hv trim5b_hv m1_23030_n25080# AGND m1_4100_n29230#
+ sky130_fd_pr__nfet_g5v0d10v5_LHNF5N
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_25 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_14 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_01v8_EPRAC4_0 Vout DVDD m1_36250_n26840# DVDD sky130_fd_pr__pfet_01v8_EPRAC4
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_33 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_22 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_11 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_01v8_HWT53N_2 DGND m1_34800_n26840# m1_36250_n26840# DGND sky130_fd_pr__nfet_01v8_HWT53N
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_26 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_15 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_LHNF5N_1 res_p_bot m1_4100_n28430# trim5b_hv trim5b_hv
+ res_p_bot trim5b_hv trim5b_hv res_p_bot AGND m1_4100_n28430# sky130_fd_pr__nfet_g5v0d10v5_LHNF5N
Xsky130_fd_pr__pfet_01v8_EPRAC4_1 m1_34800_n26840# DVDD m1_35900_10510# DVDD sky130_fd_pr__pfet_01v8_EPRAC4
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_34 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_23 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_12 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_LHNF5N_2 m1_23030_n25080# m1_4100_n28430# trim5_hv trim5_hv
+ m1_23030_n25080# trim5_hv trim5_hv m1_23030_n25080# AGND m1_4100_n28430# sky130_fd_pr__nfet_g5v0d10v5_LHNF5N
Xsky130_fd_pr__pfet_g5v0d10v5_Q8UPKT_0 m1_29940_7140# AVDD m1_29940_7140# m1_29940_7140#
+ AVDD AVDD m1_29860_5120# AVDD m1_29860_5120# AVDD m1_29940_7140# sky130_fd_pr__pfet_g5v0d10v5_Q8UPKT
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_27 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_16 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_01v8_EPRAC4_2 m1_36250_n26840# DVDD m1_34800_n26840# DVDD sky130_fd_pr__pfet_01v8_EPRAC4
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_35 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_24 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_28 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_17 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_LHNF5N_3 m1_27260_n27254# m1_23030_n25080# trim3b_hv
+ trim3b_hv m1_27260_n27254# trim3b_hv trim3b_hv m1_27260_n27254# AGND m1_23030_n25080#
+ sky130_fd_pr__nfet_g5v0d10v5_LHNF5N
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_25 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_LHNF5N_4 res_p_bot m1_4100_n29230# trim5_hv trim5_hv
+ res_p_bot trim5_hv trim5_hv res_p_bot AGND m1_4100_n29230# sky130_fd_pr__nfet_g5v0d10v5_LHNF5N
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_29 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_18 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_26 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_15 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_LHNF5N_5 res_p_bot m1_27260_n27254# trim4b_hv trim4b_hv
+ res_p_bot trim4b_hv trim4b_hv res_p_bot AGND m1_27260_n27254# sky130_fd_pr__nfet_g5v0d10v5_LHNF5N
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_19 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_27 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_16 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_MRHAE7_0 m1_30900_4740# AGND AGND m1_30900_4740# sky130_fd_pr__nfet_g5v0d10v5_MRHAE7
Xsky130_fd_pr__pfet_g5v0d10v5_X332GA_0 trim3b_hv trim3b_hv AVDD m1_33660_n22250# AVDD
+ AVDD sky130_fd_pr__pfet_g5v0d10v5_X332GA
Xsky130_fd_pr__nfet_g5v0d10v5_4RA4DJ_0 hyst1_hv AGND m1_32060_n3340# m1_32060_n3340#
+ AGND AGND m1_32060_n3340# hyst1_hv hyst1_hv AGND hyst1_hv AGND hyst1_hv hyst1_hv
+ AGND m1_32060_n3340# hyst1_hv hyst1_hv sky130_fd_pr__nfet_g5v0d10v5_4RA4DJ
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_17 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|0] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|0] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|0] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|0] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|0] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|0] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|0] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|0] res_p_bot res_p_bot casc_p casc_p AVDD
+ m1_11260_n21330# m1_11260_n21330# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|0] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|0] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|0] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|0] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|0] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|0] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|0] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|0] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|0] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|0] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|0] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|0] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|0] m1_23030_n25080# m1_23030_n25080# casc_p
+ casc_p AVDD m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|0] m1_23030_n25080# m1_23030_n25080# casc_p
+ casc_p AVDD m1_33657_n21336# m1_33657_n21336# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|0] m1_23030_n25080# m1_23030_n25080# casc_p
+ casc_p AVDD m1_33657_n21336# m1_33657_n21336# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|0] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|1] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|1] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|1] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|1] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|1] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|1] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|1] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|1] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|1] m1_12400_n19010# m1_12400_n19010# casc_p
+ casc_p AVDD m1_12860_n19530# m1_12860_n19530# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|1] m1_12400_n19010# m1_12400_n19010# casc_p
+ casc_p AVDD m1_12860_n19530# m1_12860_n19530# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|1] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|1] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|1] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|1] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|1] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|1] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|1] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|1] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|1] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|1] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|1] m1_23030_n25080# m1_23030_n25080# casc_p
+ casc_p AVDD m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|1] m1_23030_n25080# m1_23030_n25080# casc_p
+ casc_p AVDD m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|1] m1_23030_n25080# m1_23030_n25080# casc_p
+ casc_p AVDD m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|1] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|2] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|2] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|2] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|2] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|2] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|2] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|2] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|2] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|2] bias_var_n bias_var_n casc_p casc_p AVDD
+ m1_12860_n17730# m1_12860_n17730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|2] bias_var_n bias_var_n casc_p casc_p AVDD
+ m1_12860_n17730# m1_12860_n17730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|2] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|2] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|2] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|2] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|2] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|2] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|2] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|2] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|2] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|2] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|2] m1_420_n29120# m1_420_n29120# casc_p
+ casc_p AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|2] m1_420_n29120# m1_420_n29120# casc_p
+ casc_p AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|2] m1_420_n29120# m1_420_n29120# casc_p
+ casc_p AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|2] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|3] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|3] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|3] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|3] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|3] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|3] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|3] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|3] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|3] m1_2120_n22080# m1_2120_n22080# casc_p
+ casc_p AVDD m1_12860_n15930# m1_12860_n15930# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|3] m1_2120_n22080# m1_2120_n22080# casc_p
+ casc_p AVDD m1_12860_n15930# m1_12860_n15930# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|3] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|3] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|3] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|3] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|3] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|3] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|3] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|3] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|3] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|3] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|3] m1_420_n29120# m1_420_n29120# casc_p
+ casc_p AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|3] m1_420_n29120# m1_420_n29120# casc_p
+ casc_p AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|3] m1_420_n29120# m1_420_n29120# casc_p
+ casc_p AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|3] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|4] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|4] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|4] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|4] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|4] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|4] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|4] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|4] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|4] m1_2120_n22080# m1_2120_n22080# casc_p
+ casc_p AVDD m1_12860_n14130# m1_12860_n14130# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|4] m1_2120_n22080# m1_2120_n22080# casc_p
+ casc_p AVDD m1_12860_n14130# m1_12860_n14130# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|4] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|4] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|4] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|4] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|4] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|4] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|4] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|4] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|4] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|4] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|4] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|4] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|4] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|4] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|5] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|5] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|5] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|5] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|5] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|5] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|5] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|5] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|5] m1_12860_n11800# m1_12860_n11800# casc_p
+ casc_p AVDD m1_7790_4530# m1_7790_4530# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|5] m1_12860_n11800# m1_12860_n11800# casc_p
+ casc_p AVDD m1_7790_4530# m1_7790_4530# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|5] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|5] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|5] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|5] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|5] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|5] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|5] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|5] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|5] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|5] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|5] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|5] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|5] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|5] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|6] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|6] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|6] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|6] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|6] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|6] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|6] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|6] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|6] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|6] casc_p casc_p casc_p casc_p AVDD casc_p
+ casc_p sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|6] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|6] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|6] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|6] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|6] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|6] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|6] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|6] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|6] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|6] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|6] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|6] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|6] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|6] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[0|7] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[1|7] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[2|7] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[3|7] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[4|7] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[5|7] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[6|7] Vxp Vxp casc_p casc_p AVDD m1_1420_n21240#
+ m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[7|7] m1_11180_n8390# m1_11180_n8390# m1_11180_n8390#
+ m1_11180_n8390# AVDD m1_11260_n8730# m1_11260_n8730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[8|7] m1_11180_n8390# m1_11180_n8390# m1_11180_n8390#
+ m1_11180_n8390# AVDD m1_11260_n8730# m1_11260_n8730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[9|7] m1_11180_n8390# m1_11180_n8390# m1_11180_n8390#
+ m1_11180_n8390# AVDD m1_11260_n8730# m1_11260_n8730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[10|7] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[11|7] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[12|7] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[13|7] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[14|7] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[15|7] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[16|7] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[17|7] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[18|7] Vom Vom casc_p casc_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[19|7] Vop Vop casc_p casc_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[20|7] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_32060_n8730# m1_32060_n8730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[21|7] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_32060_n8730# m1_32060_n8730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[22|7] m1_31820_n13600# m1_31820_n13600# casc_p
+ casc_p AVDD m1_32060_n8730# m1_32060_n8730# sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__pfet_g5v0d10v5_GHE6BF_0[23|7] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_GHE6BF
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[0|0] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[1|0] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[2|0] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[3|0] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[4|0] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[5|0] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[6|0] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[7|0] m1_11260_n4491# AGND bias_n AGND AGND
+ m1_11260_n4491# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[8|0] m1_12840_n4260# AGND bias_n m1_12600_n4860#
+ AGND m1_12840_n4260# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[9|0] m1_14440_n4260# AGND bias_n m1_14200_n4860#
+ AGND m1_14440_n4260# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[10|0] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[11|0] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[12|0] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[13|0] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[14|0] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[15|0] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[16|0] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[17|0] m1_2500_n30560# AGND Vom AGND AGND m1_2500_n30560#
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[18|0] Vfold_bot_m AGND Vom AGND AGND Vfold_bot_m
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[19|0] m1_2500_n30560# AGND Vom AGND AGND m1_2500_n30560#
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[20|0] m1_32060_n4490# m1_32060_n3340# bias_n
+ m1_32060_n3340# AGND m1_32060_n4490# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[21|0] m1_32060_n4490# m1_32060_n3340# bias_n
+ m1_32060_n3340# AGND m1_32060_n4490# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[22|0] m1_32060_n4490# m1_32060_n3340# bias_n
+ m1_32060_n3340# AGND m1_32060_n4490# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[23|0] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[0|1] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[1|1] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[2|1] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[3|1] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[4|1] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[5|1] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[6|1] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[7|1] m1_11260_n2671# AGND bias_n AGND AGND
+ m1_11260_n2671# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[8|1] m1_12860_n2671# AGND bias_n AGND AGND
+ m1_12860_n2671# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[9|1] m1_14459_n2671# AGND bias_n AGND AGND
+ m1_14459_n2671# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[10|1] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[11|1] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[12|1] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[13|1] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[14|1] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[15|1] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[16|1] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[17|1] m1_2500_n30560# AGND Vom AGND AGND m1_2500_n30560#
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[18|1] Vfold_bot_m AGND Vom AGND AGND Vfold_bot_m
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[19|1] m1_2500_n30560# AGND Vom AGND AGND m1_2500_n30560#
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[20|1] m1_32060_n4490# m1_32060_n3340# bias_n
+ m1_32060_n3340# AGND m1_32060_n4490# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[21|1] m1_33659_n2671# m1_33660_n1540# bias_n
+ m1_33660_n1540# AGND m1_33659_n2671# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[22|1] m1_33659_n2671# AGND AGND m1_33660_n1540#
+ AGND AGND bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[23|1] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[0|2] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[1|2] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[2|2] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[3|2] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[4|2] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[5|2] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[6|2] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[7|2] bias_n AGND bias_n AGND AGND bias_n bias_n
+ sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[8|2] casc_n AGND bias_n AGND AGND casc_n bias_n
+ sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[9|2] bias_var_n AGND bias_var_n AGND AGND bias_var_n
+ bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[10|2] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[11|2] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[12|2] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[13|2] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[14|2] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[15|2] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[16|2] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[17|2] m1_2500_n30560# AGND Vom AGND AGND m1_2500_n30560#
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[18|2] Vfold_bot_m AGND Vom AGND AGND Vfold_bot_m
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[19|2] Vfold_bot_m AGND Vom AGND AGND Vfold_bot_m
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[20|2] m1_32060_n890# AGND m1_12400_n19010#
+ AGND AGND m1_32060_n890# m1_12400_n19010# sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[21|2] m1_32060_n890# AGND m1_12400_n19010#
+ AGND AGND m1_32060_n890# m1_12400_n19010# sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[22|2] m1_32060_n890# AGND m1_12400_n19010#
+ AGND AGND m1_32060_n890# m1_12400_n19010# sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[23|2] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[0|3] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[1|3] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[2|3] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[3|3] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[4|3] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[5|3] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[6|3] m1_1400_n4380# AGND bias_n AGND AGND m1_1400_n4380#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[7|3] bias_n m1_11240_2060# ibias m1_11240_2060#
+ AGND m1_11860_1120# ibias sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[8|3] m1_11860_1120# m1_12840_2060# ibias m1_12840_2060#
+ AGND ibias ibias sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[9|3] m1_12400_n19010# AGND m1_12400_n19010#
+ AGND AGND m1_12400_n19010# m1_12400_n19010# sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[10|3] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[11|3] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[12|3] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[13|3] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[14|3] Vfold_bot_m AGND bias_var_n AGND AGND
+ Vfold_bot_m bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[15|3] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[16|3] m1_2500_n30560# AGND bias_var_n AGND
+ AGND m1_2500_n30560# bias_var_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[17|3] m1_2500_n30560# AGND Vom AGND AGND m1_2500_n30560#
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[18|3] Vfold_bot_m AGND Vom AGND AGND Vfold_bot_m
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[19|3] Vfold_bot_m AGND Vom AGND AGND Vfold_bot_m
+ Vom sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[20|3] m1_32060_910# m1_32060_2060# bias_n m1_32060_2060#
+ AGND m1_32060_910# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[21|3] m1_32060_910# m1_32060_2060# bias_n m1_32060_2060#
+ AGND m1_32060_910# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[22|3] m1_35259_929# m1_35270_2060# bias_n m1_35270_2060#
+ AGND m1_35259_929# bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_WGHV7X_0[23|3] m1_36870_930# AGND bias_n AGND AGND m1_37480_930#
+ bias_n sky130_fd_pr__nfet_g5v0d10v5_WGHV7X
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_28 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_MRHAE7_1 DGND DGND m1_35900_10510# m1_30900_4740# sky130_fd_pr__nfet_g5v0d10v5_MRHAE7
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_29 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_18 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_0 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_19 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_1 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_2 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_0 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_3 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_1 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_2 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_4 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_LURNA9_0 m1_32060_n4840# m1_2500_5340# m1_32060_n4840#
+ m1_34800_n26840# m1_34800_n26840# m1_32060_n4840# AGND m1_2500_5340# m1_34800_n26840#
+ m1_34800_n26840# m1_2500_5340# m1_34800_n26840# m1_2500_5340# m1_2500_5340# m1_34800_n26840#
+ m1_34800_n26840# m1_34800_n26840# m1_32060_n4840# sky130_fd_pr__nfet_g5v0d10v5_LURNA9
Xsky130_fd_pr__nfet_g5v0d10v5_RM8L2M_0 AGND m1_29880_4800# m1_30900_4740# AGND sky130_fd_pr__nfet_g5v0d10v5_RM8L2M
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_3 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_N8ANR9_0 m1_23040_4590# m1_4100_9160# m1_23040_4590#
+ AVDD level_shifter_up_7/xb_hv level_shifter_up_7/xb_hv level_shifter_up_7/xb_hv
+ level_shifter_up_7/xb_hv m1_23040_4590# m1_4100_9160# sky130_fd_pr__pfet_g5v0d10v5_N8ANR9
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_5 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__nfet_g5v0d10v5_LURNA9_1 m1_32060_n4840# m1_2500_6140# m1_32060_n4840#
+ m1_36250_n26840# m1_36250_n26840# m1_32060_n4840# AGND m1_2500_6140# m1_36250_n26840#
+ m1_36250_n26840# m1_2500_6140# m1_36250_n26840# m1_2500_6140# m1_2500_6140# m1_36250_n26840#
+ m1_36250_n26840# m1_36250_n26840# m1_32060_n4840# sky130_fd_pr__nfet_g5v0d10v5_LURNA9
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[0|0] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[1|0] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[2|0] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[3|0] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[4|0] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[5|0] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[6|0] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[7|0] casc_n casc_n casc_p casc_p m1_11260_n4491#
+ AGND m1_11260_n4491# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[8|0] casc_n casc_n m1_11180_n8390# m1_12600_n4860#
+ m1_12850_n4460# AGND m1_12850_n4460# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[9|0] casc_n casc_n m1_12860_n11800# m1_14200_n4860#
+ m1_14450_n4460# AGND m1_14450_n4460# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[10|0] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[11|0] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[12|0] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[13|0] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[14|0] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[15|0] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[16|0] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[17|0] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[18|0] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[19|0] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[20|0] casc_n casc_n m1_32060_n4840# m1_32060_n4840#
+ m1_32060_n4490# AGND m1_32060_n4490# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[21|0] casc_n casc_n m1_32060_n4840# m1_32060_n4840#
+ m1_32060_n4490# AGND m1_32060_n4490# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[22|0] casc_n casc_n m1_32060_n4840# m1_32060_n4840#
+ m1_32060_n4490# AGND m1_32060_n4490# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[23|0] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[0|1] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[1|1] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[2|1] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[3|1] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[4|1] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[5|1] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[6|1] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[7|1] casc_n casc_n bias_p bias_p m1_11260_n2671#
+ AGND m1_11260_n2671# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[8|1] casc_n casc_n m1_9080_4100# m1_9080_4100#
+ m1_12860_n2671# AGND m1_12860_n2671# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[9|1] casc_n casc_n m1_2120_n22080# m1_2120_n22080#
+ m1_14459_n2671# AGND m1_14459_n2671# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[10|1] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[11|1] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[12|1] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[13|1] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[14|1] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[15|1] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[16|1] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[17|1] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[18|1] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[19|1] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[20|1] casc_n casc_n m1_32060_n4840# m1_32060_n4840#
+ m1_32060_n4490# AGND m1_32060_n4490# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[21|1] casc_n casc_n m1_32060_n4840# m1_32060_n4840#
+ m1_33659_n2671# AGND m1_33659_n2671# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[22|1] casc_n casc_n casc_n m1_32060_n4840#
+ m1_33659_n2671# AGND casc_n sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[23|1] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[0|2] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[1|2] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[2|2] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[3|2] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[4|2] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[5|2] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[6|2] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[7|2] casc_n casc_n casc_n casc_n casc_n AGND
+ casc_n sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[8|2] ibias ibias AVDD AVDD casc_n AGND casc_n
+ sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[9|2] casc_n casc_n casc_n casc_n casc_n AGND
+ casc_n sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[10|2] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[11|2] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[12|2] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[13|2] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[14|2] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[15|2] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[16|2] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[17|2] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[18|2] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[19|2] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[20|2] casc_n casc_n m1_420_6500# m1_420_6500#
+ m1_32060_n890# AGND m1_32060_n890# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[21|2] casc_n casc_n m1_420_6500# m1_420_6500#
+ m1_32060_n890# AGND m1_32060_n890# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[22|2] casc_n casc_n m1_420_6500# m1_420_6500#
+ m1_32060_n890# AGND m1_32060_n890# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[23|2] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[0|3] AGND AGND AGND AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[1|3] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[2|3] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[3|3] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[4|3] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[5|3] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[6|3] casc_n casc_n Vxm Vxm m1_1400_n4380# AGND
+ m1_1400_n4380# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[7|3] casc_n casc_n casc_n casc_n casc_n AGND
+ casc_n sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[8|3] casc_n casc_n casc_n casc_n casc_n AGND
+ casc_n sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[9|3] casc_n casc_n casc_n casc_n casc_n AGND
+ casc_n sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[10|3] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[11|3] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[12|3] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[13|3] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[14|3] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[15|3] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[16|3] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[17|3] casc_n casc_n Vop Vop m1_2500_n30560#
+ AGND m1_2500_n30560# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[18|3] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[19|3] casc_n casc_n Vom Vom Vfold_bot_m AGND
+ Vfold_bot_m sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[20|3] casc_n casc_n m1_23040_4590# m1_23040_4590#
+ m1_32060_910# AGND m1_32060_910# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[21|3] casc_n casc_n m1_23040_4590# m1_23040_4590#
+ m1_32060_910# AGND m1_32060_910# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[22|3] casc_n casc_n m1_23040_4590# m1_23040_4590#
+ m1_35259_929# AGND m1_35259_929# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__nfet_g5v0d10v5_CDNABP_0[23|3] casc_n casc_n m1_29940_7140# m1_25710_11400#
+ m1_36870_930# AGND m1_37480_930# sky130_fd_pr__nfet_g5v0d10v5_CDNABP
Xsky130_fd_pr__pfet_g5v0d10v5_N8ANR9_1 m1_25710_11400# m1_27260_9746# m1_25710_11400#
+ AVDD level_shifter_up_6/x_hv level_shifter_up_6/x_hv level_shifter_up_6/x_hv level_shifter_up_6/x_hv
+ m1_25710_11400# m1_27260_9746# sky130_fd_pr__pfet_g5v0d10v5_N8ANR9
Xsky130_fd_pr__pfet_g5v0d10v5_6UJQA2_0 AVDD bias_p AVDD bias_p AVDD en_hv en_hv en_hv
+ en_hv bias_p sky130_fd_pr__pfet_g5v0d10v5_6UJQA2
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_6 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_4 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_5 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_N8ANR9_2 m1_27260_9746# m1_23040_4590# m1_27260_9746#
+ AVDD level_shifter_up_8/x_hv level_shifter_up_8/x_hv level_shifter_up_8/x_hv level_shifter_up_8/x_hv
+ m1_27260_9746# m1_23040_4590# sky130_fd_pr__pfet_g5v0d10v5_N8ANR9
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|0] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|0] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|0] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|0] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|0] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|0] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|0] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|0] bias_p AVDD AVDD bias_p AVDD m1_11260_n21330#
+ m1_11260_n21330# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|0] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|0] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|0] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|0] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|0] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|0] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|0] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|0] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|0] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|0] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|0] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|0] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|0] bias_p m1_32060_n22250# AVDD bias_p m1_32060_n22250#
+ m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|0] bias_p m1_33660_n22250# AVDD bias_p m1_33660_n22250#
+ m1_33657_n21336# m1_33657_n21336# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|0] bias_p m1_33660_n22250# AVDD bias_p m1_33660_n22250#
+ m1_33657_n21336# m1_33657_n21336# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|0] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|1] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|1] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|1] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|1] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|1] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|1] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|1] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|1] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_12860_n19530# m1_12860_n19530# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_12860_n19530# m1_12860_n19530# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|1] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|1] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|1] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|1] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|1] bias_p m1_32060_n22250# AVDD bias_p m1_32060_n22250#
+ m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|1] bias_p m1_32060_n22250# AVDD bias_p m1_32060_n22250#
+ m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|1] bias_p m1_32060_n22250# AVDD bias_p m1_32060_n22250#
+ m1_31740_n21330# m1_31740_n21330# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|1] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|2] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|2] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_12860_n17730# m1_12860_n17730# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_12860_n17730# m1_12860_n17730# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|2] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|2] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|2] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|2] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|2] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|2] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|2] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|2] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|2] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|2] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|2] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|2] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|3] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|3] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_12860_n15930# m1_12860_n15930# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_12860_n15930# m1_12860_n15930# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|3] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|3] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|3] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|3] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|3] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|3] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|3] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|3] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|3] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|3] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|3] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_31580_n17650# m1_31580_n17650# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|3] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|4] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|4] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|4] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|4] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|4] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|4] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|4] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|4] bias_p AVDD AVDD bias_p AVDD m1_11260_n14130#
+ m1_11260_n14130# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_12860_n14130# m1_12860_n14130# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_12860_n14130# m1_12860_n14130# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|4] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|4] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|4] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|4] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|4] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|4] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|4] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|4] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|5] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|5] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|5] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|5] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|5] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|5] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|5] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|5] bias_p m1_11260_n14130# AVDD bias_p m1_11260_n14130#
+ m1_7790_4530# m1_7790_4530# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_7790_4530# m1_7790_4530# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_7790_4530# m1_7790_4530# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|5] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|5] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|5] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|5] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|5] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|5] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|5] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|5] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|6] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|6] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|6] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|6] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|6] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|6] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|6] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|6] bias_p AVDD AVDD bias_p AVDD bias_p bias_p
+ sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|6] bias_p AVDD AVDD bias_p AVDD bias_p bias_p
+ sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|6] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|6] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|6] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|6] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|6] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|6] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|6] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|6] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|6] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|6] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|6] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|6] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|6] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|6] bias_p m1_32060_n15040# AVDD bias_p m1_32060_n15040#
+ m1_31600_n14050# m1_31600_n14050# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|6] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[0|7] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[1|7] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[2|7] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[3|7] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[4|7] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[5|7] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[6|7] m1_2120_n22080# AVDD AVDD m1_2120_n22080#
+ AVDD m1_1420_n21240# m1_1420_n21240# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[7|7] m1_11180_n8390# AVDD AVDD m1_11180_n8390#
+ AVDD m1_11260_n8730# m1_11260_n8730# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[8|7] casc_p m1_11260_n8730# AVDD casc_p m1_11260_n8730#
+ casc_p casc_p sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[9|7] casc_p m1_11260_n8730# AVDD casc_p m1_11260_n8730#
+ casc_p casc_p sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[10|7] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[11|7] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[12|7] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[13|7] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[14|7] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[15|7] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_6140# m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[16|7] m1_12860_n11800# AVDD AVDD m1_12860_n11800#
+ AVDD m1_2500_5340# m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[17|7] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[18|7] bias_p AVDD AVDD bias_p AVDD m1_2500_5340#
+ m1_2500_5340# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[19|7] bias_p AVDD AVDD bias_p AVDD m1_2500_6140#
+ m1_2500_6140# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[20|7] bias_p m1_32060_n9640# AVDD bias_p m1_32060_n9640#
+ m1_32060_n8730# m1_32060_n8730# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[21|7] bias_p m1_32060_n9640# AVDD bias_p m1_32060_n9640#
+ m1_32060_n8730# m1_32060_n8730# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[22|7] bias_p m1_32060_n9640# AVDD bias_p m1_32060_n9640#
+ m1_32060_n8730# m1_32060_n8730# sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__pfet_g5v0d10v5_CS979Q_0[23|7] AVDD AVDD AVDD AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_CS979Q
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_7 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_2CKAKF_0 m1_32060_n15040# AVDD AVDD m1_32060_n15040#
+ hyst1b_hv hyst1b_hv hyst1b_hv m1_32060_n15040# m1_32060_n15040# AVDD hyst1b_hv hyst1b_hv
+ hyst1b_hv hyst1b_hv AVDD AVDD hyst1b_hv hyst1b_hv hyst1b_hv AVDD hyst1b_hv hyst1b_hv
+ m1_32060_n15040# hyst1b_hv hyst1b_hv m1_32060_n15040# hyst1b_hv AVDD AVDD hyst1b_hv
+ AVDD m1_32060_n15040# AVDD m1_32060_n15040# sky130_fd_pr__pfet_g5v0d10v5_2CKAKF
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_8 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_6 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_N8ANR9_3 m1_25710_11400# m1_4100_9160# m1_25710_11400#
+ AVDD level_shifter_up_7/x_hv level_shifter_up_7/x_hv level_shifter_up_7/x_hv level_shifter_up_7/x_hv
+ m1_25710_11400# m1_4100_9160# sky130_fd_pr__pfet_g5v0d10v5_N8ANR9
Xsky130_fd_pr__nfet_g5v0d10v5_EEFBWQ_0 AGND AGND res_p_bot res_p_bot sky130_fd_pr__nfet_g5v0d10v5_EEFBWQ
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_7 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_N8ANR9_4 m1_25710_11400# m1_4100_8360# m1_25710_11400#
+ AVDD level_shifter_up_7/xb_hv level_shifter_up_7/xb_hv level_shifter_up_7/xb_hv
+ level_shifter_up_7/xb_hv m1_25710_11400# m1_4100_8360# sky130_fd_pr__pfet_g5v0d10v5_N8ANR9
Xsky130_fd_pr__nfet_g5v0d10v5_T8W2FW_9 AGND AGND AGND AGND sky130_fd_pr__nfet_g5v0d10v5_T8W2FW
Xlevel_shifter_up_0 AVDD trim[5] trim5_hv trim5b_hv DVDD DGND m1_33128_n32592# AGND
+ level_shifter_up
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_8 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xsky130_fd_pr__pfet_g5v0d10v5_N8ANR9_5 m1_23040_4590# m1_4100_8360# m1_23040_4590#
+ AVDD level_shifter_up_7/x_hv level_shifter_up_7/x_hv level_shifter_up_7/x_hv level_shifter_up_7/x_hv
+ m1_23040_4590# m1_4100_8360# sky130_fd_pr__pfet_g5v0d10v5_N8ANR9
Xsky130_fd_pr__pfet_g5v0d10v5_9432CF_0 AVDD hyst0b_hv hyst0b_hv AVDD hyst0b_hv m1_32060_n9640#
+ m1_32060_n9640# hyst0b_hv hyst0b_hv AVDD hyst0b_hv m1_32060_n9640# AVDD m1_32060_n9640#
+ sky130_fd_pr__pfet_g5v0d10v5_9432CF
Xlevel_shifter_up_1 AVDD hyst[0] hyst0_hv hyst0b_hv DVDD DGND m1_38128_n32592# AGND
+ level_shifter_up
Xsky130_fd_pr__pfet_g5v0d10v5_PNRDLC_9 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_g5v0d10v5_PNRDLC
Xlevel_shifter_up_2 AVDD hyst[1] hyst1_hv hyst1b_hv DVDD DGND m1_37128_n32592# AGND
+ level_shifter_up
Xsky130_fd_pr__nfet_g5v0d10v5_M7X63G_81 Vxm m1_2500_5340# Vinp AGND sky130_fd_pr__nfet_g5v0d10v5_M7X63G
Xsky130_fd_pr__pfet_g5v0d10v5_REE66T_0 m1_34800_n26840# Vfold_bot_m Vfold_bot_m m1_34800_n26840#
+ m1_31820_n13600# m1_34800_n26840# m1_31820_n13600# Vfold_bot_m m1_34800_n26840#
+ m1_34800_n26840# m1_31820_n13600# m1_34800_n26840# m1_34800_n26840# m1_34800_n26840#
+ m1_31820_n13600# Vfold_bot_m AVDD Vfold_bot_m sky130_fd_pr__pfet_g5v0d10v5_REE66T
Xsky130_fd_pr__pfet_g5v0d10v5_2432J2_1 AVDD trim4b_hv trim4b_hv trim4b_hv m1_32060_n22250#
+ trim4b_hv AVDD AVDD m1_32060_n22250# AVDD sky130_fd_pr__pfet_g5v0d10v5_2432J2
.ends

.subckt sky130_fd_pr__nfet_01v8_PVEW3M a_n210_n274# a_50_n100# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n210_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_XPB8Y6 a_n50_n297# a_50_n200# a_n108_n200# w_n246_n419#
X0 a_50_n200# a_n50_n297# a_n108_n200# w_n246_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt Stage0_clk_inv dvddb clka clk clkb dvss
XXM6 dvss clkb dvss clk sky130_fd_pr__nfet_01v8_PVEW3M
XXM8 clkb clka dvddb dvddb sky130_fd_pr__pfet_01v8_XPB8Y6
XXM21 dvss clka dvss clkb sky130_fd_pr__nfet_01v8_PVEW3M
XXM22 clk clkb dvddb dvddb sky130_fd_pr__pfet_01v8_XPB8Y6
.ends

.subckt sky130_fd_pr__pfet_01v8_hvt_3HBZVM a_n158_n300# w_n296_n519# a_n100_n397#
+ a_100_n300#
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n296_n519# sky130_fd_pr__pfet_01v8_hvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_WSEQJ8 a_50_n200# a_n242_n422# a_n108_n200# a_n50_n288#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n242_n422# sky130_fd_pr__nfet_03v3_nvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_3HY9VM w_n296_n419# a_n100_n297# a_100_n200# a_n158_n200#
X0 a_100_n200# a_n100_n297# a_n158_n200# w_n296_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_UNEQ2N a_n252_n322# a_50_n100# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n252_n322# sky130_fd_pr__nfet_03v3_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt Stage2_latch dvdd enab clkb vout oneg opos dvss dvddb
XXM12 dvddb dvddb clkb m1_683_n2348# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM15 dvss dvss m2_1568_n2406# clkb sky130_fd_pr__nfet_03v3_nvt_WSEQJ8
XXM18 dvss dvss vout m1_683_n2348# sky130_fd_pr__nfet_01v8_PVEW3M
XXM19 dvddb m1_683_n2348# dvddb vout sky130_fd_pr__pfet_01v8_3HY9VM
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_0 dvddb dvddb clkb m2_1331_n391# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM1 dvddb dvddb m2_1331_n391# m1_683_n2348# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_1 dvddb dvddb m1_683_n2348# m2_1331_n391# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_3 dvddb dvddb m1_683_n2348# m2_1331_n391# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_2 dvddb dvddb clkb m2_1331_n391# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM2 dvss m1_1866_n2368# m1_683_n2348# opos sky130_fd_pr__nfet_03v3_nvt_UNEQ2N
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_4 dvdd dvdd enab dvddb sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM3 dvss m2_1568_n2406# m1_1866_n2368# m2_1331_n391# sky130_fd_pr__nfet_03v3_nvt_UNEQ2N
Xsky130_fd_pr__pfet_01v8_hvt_3HBZVM_5 dvdd dvdd enab dvddb sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM4 dvss m1_2747_n2368# m2_1331_n391# oneg sky130_fd_pr__nfet_03v3_nvt_UNEQ2N
XXM5 dvss m2_1568_n2406# m1_2747_n2368# m1_683_n2348# sky130_fd_pr__nfet_03v3_nvt_UNEQ2N
XXM10 dvddb dvddb clkb m1_683_n2348# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
XXM11 dvddb dvddb m2_1331_n391# m1_683_n2348# sky130_fd_pr__pfet_01v8_hvt_3HBZVM
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_FGL9FS a_29_n597# a_n287_n500# a_n229_n597# a_287_n597#
+ a_229_n500# w_n745_n797# a_n545_n500# a_n487_n597# a_n29_n500# a_487_n500#
X0 a_487_n500# a_287_n597# a_229_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X1 a_229_n500# a_29_n597# a_n29_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_n29_n500# a_n229_n597# a_n287_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_n287_n500# a_n487_n597# a_n545_n500# w_n745_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_E2TVSU a_1261_n500# a_n1319_n500# a_29_n597#
+ a_n287_n500# a_n1061_n500# a_n745_n597# a_803_n597# a_745_n500# a_n229_n597# a_287_n597#
+ a_n1003_n597# a_229_n500# w_n1519_n797# a_n545_n500# a_1061_n597# a_1003_n500# a_n487_n597#
+ a_n1261_n597# a_n29_n500# a_545_n597# a_487_n500# a_n803_n500#
X0 a_n1061_n500# a_n1261_n597# a_n1319_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X1 a_1003_n500# a_803_n597# a_745_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X2 a_487_n500# a_287_n597# a_229_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X3 a_745_n500# a_545_n597# a_487_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X4 a_1261_n500# a_1061_n597# a_1003_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X5 a_229_n500# a_29_n597# a_n29_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X6 a_n29_n500# a_n229_n597# a_n287_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X7 a_n545_n500# a_n745_n597# a_n803_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X8 a_n287_n500# a_n487_n597# a_n545_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X9 a_n803_n500# a_n1003_n597# a_n1061_n500# w_n1519_n797# sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y a_50_n500# a_n242_n722# a_n108_n500# a_n50_n588#
X0 a_50_n500# a_n50_n588# a_n108_n500# a_n242_n722# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y a_50_n500# a_n242_n722# a_n108_n500# a_n50_n588#
X0 a_50_n500# a_n50_n588# a_n108_n500# a_n242_n722# sky130_fd_pr__nfet_03v3_nvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.5
.ends

.subckt Stage1 avdd clka vinn vinp oneg opos avss dvdd dvss w_608_n4573# enab
Xx1 clka dvdd dvss avdd avdd x1/X avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xx2 enab dvdd dvss avdd avdd x2/X avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
XXM3_2 vinp oneg vinp vinp oneg li_n3_908# li_n3_908# vinp li_n3_908# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_FGL9FS
XXM1_1 avdd avdd x2/X avdd li_1882_n1884# x2/X x2/X avdd x2/X x2/X x2/X avdd avdd
+ li_1882_n1884# x2/X li_1882_n1884# x2/X x2/X li_1882_n1884# x2/X li_1882_n1884#
+ avdd sky130_fd_pr__pfet_g5v0d10v5_E2TVSU
XXM1_2 avdd avdd x2/X avdd li_1882_n1884# x2/X x2/X avdd x2/X x2/X x2/X avdd avdd
+ li_1882_n1884# x2/X li_1882_n1884# x2/X x2/X li_1882_n1884# x2/X li_1882_n1884#
+ avdd sky130_fd_pr__pfet_g5v0d10v5_E2TVSU
XXM5 opos w_608_n4573# w_608_n4573# x1/X sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y
XXM6_1 li_n3_908# li_n3_908# x1/X li_n3_908# li_1882_n1884# x1/X x1/X li_n3_908# x1/X
+ x1/X x1/X li_n3_908# li_1882_n1884# li_1882_n1884# x1/X li_1882_n1884# x1/X x1/X
+ li_1882_n1884# x1/X li_1882_n1884# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_E2TVSU
XXM6_2 li_n3_908# li_n3_908# x1/X li_n3_908# li_1882_n1884# x1/X x1/X li_n3_908# x1/X
+ x1/X x1/X li_n3_908# li_1882_n1884# li_1882_n1884# x1/X li_1882_n1884# x1/X x1/X
+ li_1882_n1884# x1/X li_1882_n1884# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_E2TVSU
XXM8 oneg w_608_n4573# w_608_n4573# x1/X sky130_fd_pr__nfet_g5v0d10v5_FJGQ2Y
XXM4_2 avss avss w_608_n4573# w_608_n4573# sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y
Xsky130_fd_pr__pfet_g5v0d10v5_FGL9FS_0 vinp oneg vinp vinp oneg li_n3_908# li_n3_908#
+ vinp li_n3_908# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_FGL9FS
Xsky130_fd_pr__pfet_g5v0d10v5_FGL9FS_1 vinn opos vinn vinn opos li_n3_908# li_n3_908#
+ vinn li_n3_908# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_FGL9FS
XXM2_2 vinn opos vinn vinn opos li_n3_908# li_n3_908# vinn li_n3_908# li_n3_908# sky130_fd_pr__pfet_g5v0d10v5_FGL9FS
Xsky130_fd_pr__nfet_03v3_nvt_FJGQ2Y_0 avss avss w_608_n4573# w_608_n4573# sky130_fd_pr__nfet_03v3_nvt_FJGQ2Y
.ends

.subckt Stage0_ena_inv dvdd ena enab dvss
XXM24 dvss enab dvss ena sky130_fd_pr__nfet_01v8_PVEW3M
XXM25 ena enab dvdd dvdd sky130_fd_pr__pfet_01v8_XPB8Y6
.ends

.subckt sky130_icrg_ip__ulpcomp2 avdd ena vout vinn vinp dvss clk dvdd avss w_288_n7621#
Xx1 x3/dvddb x2/clka clk x3/clkb dvss Stage0_clk_inv
Xx3 dvdd x4/enab x3/clkb vout x3/oneg x3/opos dvss x3/dvddb Stage2_latch
Xx2 avdd x2/clka vinn vinp x3/oneg x3/opos avss dvdd dvss w_288_n7621# x4/enab Stage1
Xx4 dvdd ena x4/enab dvss Stage0_ena_inv
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLHCT5 a_n345_n200# a_29_n297# a_n129_n297# a_187_n297#
+ a_129_n200# a_n287_n297# a_287_n200# a_n29_n200# a_n187_n200# w_n545_n497#
X0 a_n187_n200# a_n287_n297# a_n345_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X1 a_287_n200# a_187_n297# a_129_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2 a_129_n200# a_29_n297# a_n29_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X3 a_n29_n200# a_n129_n297# a_n187_n200# w_n545_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KL97Y6 a_29_n297# a_n129_n297# a_129_n200# a_n29_n200#
+ w_n387_n497# a_n187_n200#
X0 a_129_n200# a_29_n297# a_n29_n200# w_n387_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X1 a_n29_n200# a_n129_n297# a_n187_n200# w_n387_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EJGQFX a_129_n200# a_29_n288# a_n129_n288# a_n321_n422#
+ a_n29_n200# a_n187_n200#
X0 a_129_n200# a_29_n288# a_n29_n200# a_n321_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X1 a_n29_n200# a_n129_n288# a_n187_n200# a_n321_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8 a_50_n200# a_n242_n422# a_n108_n200# a_n50_n288#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n242_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt simple_analog_switch on off out in vdd vss
XXM12 out off off off in off out out in vdd sky130_fd_pr__pfet_g5v0d10v5_KLHCT5
XXM14 on on out out vdd out sky130_fd_pr__pfet_g5v0d10v5_KL97Y6
XXM16 on on in in vdd in sky130_fd_pr__pfet_g5v0d10v5_KL97Y6
XXM1 out on on vss in out sky130_fd_pr__nfet_g5v0d10v5_EJGQFX
XXM3 out vss out off sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8
XXM5 in vss in off sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8
.ends

.subckt EF_SW_RST VP2 VP1 AVDD DVDD AVSS HOLD DVSS HOLDB VIN m3_2464_n194# m3_1864_n2876#
Xsimple_analog_switch_0 HOLDB HOLD VP2 VIN AVDD AVSS simple_analog_switch
Xsimple_analog_switch_1 HOLDB HOLD VIN VP1 AVDD AVSS simple_analog_switch
.ends

.subckt sky130_fd_sc_hvl__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0 ps=0 w=0.75 l=1
X2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0 ps=0 w=1 l=1
X3 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0 ps=0 w=0.75 l=1
.ends

.subckt sky130_fd_sc_hvl__nor2_1 A B VGND VNB VPB VPWR Y
X0 a_251_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.1575 pd=1.71 as=0.4275 ps=3.57 w=1.5 l=0.5
X1 Y B a_251_443# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.4275 pd=3.57 as=0.1575 ps=1.71 w=1.5 l=0.5
X2 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21375 ps=2.07 w=0.75 l=0.5
X3 VGND B Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.21375 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt EF_AMUX21x vdd1p8 a sel selcm cm vss vo vdd3p3 b dvss
Xsimple_analog_switch_2_0 sky130_fd_sc_hvl__inv_2_3/A vdd3p3 vss sky130_fd_sc_hvl__inv_2_3/Y
+ vo a simple_analog_switch_2
Xsimple_analog_switch_2_1 sky130_fd_sc_hvl__inv_2_0/A vdd3p3 vss sky130_fd_sc_hvl__inv_2_0/Y
+ vo b simple_analog_switch_2
Xsimple_analog_switch_2_2 sky130_fd_sc_hvl__inv_2_5/Y vdd3p3 vss sky130_fd_sc_hvl__inv_2_5/A
+ vo cm simple_analog_switch_2
Xsky130_fd_sc_hvl__inv_2_0 sky130_fd_sc_hvl__inv_2_0/A dvss dvss vdd3p3 vdd3p3 sky130_fd_sc_hvl__inv_2_0/Y
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_1 selcm dvss dvss vdd3p3 vdd3p3 sky130_fd_sc_hvl__inv_2_5/A
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_2 sel dvss dvss vdd3p3 vdd3p3 sky130_fd_sc_hvl__inv_2_2/Y
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_3 sky130_fd_sc_hvl__inv_2_3/A dvss dvss vdd3p3 vdd3p3 sky130_fd_sc_hvl__inv_2_3/Y
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_5 sky130_fd_sc_hvl__inv_2_5/A dvss dvss vdd3p3 vdd3p3 sky130_fd_sc_hvl__inv_2_5/Y
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__decap_8_0 dvss dvss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_8
Xsky130_fd_sc_hvl__decap_8_1 dvss dvss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_8
Xsky130_fd_sc_hvl__decap_8_2 dvss dvss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_8
Xsky130_fd_sc_hvl__decap_8_3 dvss dvss vdd3p3 vdd3p3 sky130_fd_sc_hvl__decap_8
Xsky130_fd_sc_hvl__nor2_1_0 selcm sky130_fd_sc_hvl__inv_2_2/Y dvss dvss vdd3p3 vdd3p3
+ sky130_fd_sc_hvl__inv_2_0/A sky130_fd_sc_hvl__nor2_1
Xsky130_fd_sc_hvl__nor2_1_1 sel selcm dvss dvss vdd3p3 vdd3p3 sky130_fd_sc_hvl__inv_2_3/A
+ sky130_fd_sc_hvl__nor2_1
.ends

.subckt EF_AMUX0201_ARRAY1 SELD2 SELD3 SELD0 SELD1 SELD4 D1 SELD5 SELD9 SELD8 D5 SELD7
+ D9 SELD6 D8 D7 DVSS SELD10 SELD11 VCM D11 D0 x9/selcm D4 D2 x4/selcm D10 VH DVDD
+ D6 D3 VDD VL VSS
Xx1 DVDD VH SELD3 x4/selcm VCM VSS D3 VDD VL DVSS EF_AMUX21x
Xx3 DVDD VH SELD8 x4/selcm VCM VSS D8 VDD VL DVSS EF_AMUX21x
Xx2 DVDD VH SELD4 x9/selcm VCM VSS D4 VDD VL DVSS EF_AMUX21x
Xx4 DVDD VH SELD6 x4/selcm VCM VSS D6 VDD VL DVSS EF_AMUX21x
Xx5 DVDD VH SELD0 x9/selcm VCM VSS D0 VDD VL DVSS EF_AMUX21x
Xx8 DVDD VH SELD2 x9/selcm VCM VSS D2 VDD VL DVSS EF_AMUX21x
Xx9 DVDD VH SELD11 x9/selcm VCM VSS D11 VDD VL DVSS EF_AMUX21x
Xx10 DVDD VH SELD5 x4/selcm VCM VSS D5 VDD VL DVSS EF_AMUX21x
Xx11 DVDD VH SELD1 x4/selcm VCM VSS D1 VDD VL DVSS EF_AMUX21x
Xx12 DVDD VH SELD10 x4/selcm VCM VSS D10 VDD VL DVSS EF_AMUX21x
XEF_AMUX21x_0 DVDD VH SELD9 x9/selcm VCM VSS D9 VDD VL DVSS EF_AMUX21x
XEF_AMUX21x_1 DVDD VH SELD7 x9/selcm VCM VSS D7 VDD VL DVSS EF_AMUX21x
.ends

.subckt cdac_unit_cap m3_80891_n32882# c1_81071_n33152# c2_81071_n33152#
X0 c1_81071_n33152# m3_80891_n32882# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X1 c2_81071_n33152# c1_81071_n33152# sky130_fd_pr__cap_mim_m3_2 l=7 w=7
.ends

.subckt cap_array_half cdac_unit_cap_1[4|9]/c2_81071_n33152# cdac_unit_cap_1[3|0]/m3_80891_n32882#
+ cdac_unit_cap_1[7|7]/m3_80891_n32882# cdac_unit_cap_1[6|7]/m3_80891_n32882# cdac_unit_cap_1[6|9]/m3_80891_n32882#
+ cdac_unit_cap_1[6|0]/c2_81071_n33152# cdac_unit_cap_1[2|7]/m3_80891_n32882# cdac_unit_cap_1[8|0]/m3_80891_n32882#
+ cdac_unit_cap_1[5|1]/m3_80891_n32882# cdac_unit_cap_1[3|9]/c2_81071_n33152# cdac_unit_cap_1[2|0]/m3_80891_n32882#
+ cdac_unit_cap_1[7|5]/m3_80891_n32882# cdac_unit_cap_1[5|9]/m3_80891_n32882# cdac_unit_cap_1[5|0]/c2_81071_n33152#
+ cdac_unit_cap_1[8|9]/c2_81071_n33152# cdac_unit_cap_1[4|4]/m3_80891_n32882# cdac_unit_cap_1[7|0]/m3_80891_n32882#
+ cdac_unit_cap_1[2|6]/m3_80891_n32882# cdac_unit_cap_1[2|9]/c2_81071_n33152# cdac_unit_cap_1[2|8]/m3_80891_n32882#
+ cdac_unit_cap_1[1|0]/m3_80891_n32882# cdac_unit_cap_1[4|9]/m3_80891_n32882# cdac_unit_cap_1[4|0]/c2_81071_n33152#
+ cdac_unit_cap_1[7|9]/c2_81071_n33152# cdac_unit_cap_1[6|0]/m3_80891_n32882# cdac_unit_cap_1[3|7]/m3_80891_n32882#
+ cdac_unit_cap_1[4|4]/c1_81071_n33152# cdac_unit_cap_1[1|9]/c2_81071_n33152# cdac_unit_cap_1[8|8]/m3_80891_n32882#
+ cdac_unit_cap_1[5|7]/m3_80891_n32882# cdac_unit_cap_1[1|7]/m3_80891_n32882# cdac_unit_cap_1[3|9]/m3_80891_n32882#
+ cdac_unit_cap_1[3|0]/c2_81071_n33152# cdac_unit_cap_1[5|5]/m3_80891_n32882# cdac_unit_cap_1[6|9]/c2_81071_n33152#
+ cdac_unit_cap_1[6|8]/m3_80891_n32882# cdac_unit_cap_1[8|7]/m3_80891_n32882# cdac_unit_cap_1[5|0]/m3_80891_n32882#
+ cdac_unit_cap_1[8|9]/m3_80891_n32882# cdac_unit_cap_1[8|0]/c2_81071_n33152# cdac_unit_cap_1[2|9]/m3_80891_n32882#
+ cdac_unit_cap_1[2|0]/c2_81071_n33152# cdac_unit_cap_1[5|9]/c2_81071_n33152# caparray_connect_none_8/m3_85388_n19067#
+ cdac_unit_cap_1[4|8]/m3_80891_n32882# cdac_unit_cap_1[4|0]/m3_80891_n32882# cdac_unit_cap_1[7|9]/m3_80891_n32882#
+ cdac_unit_cap_1[7|0]/c2_81071_n33152# cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_99908_n7967#
+ m4_81638_n9537# cdac_unit_cap_1[1|9]/m3_80891_n32882# cdac_unit_cap_1[1|0]/c2_81071_n33152#
+ cdac_unit_cap_1[4|7]/m3_80891_n32882#
Xcdac_unit_cap_1[0|0] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|0] cdac_unit_cap_1[1|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[1|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|0] cdac_unit_cap_1[2|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[2|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|0] cdac_unit_cap_1[3|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[3|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|0] cdac_unit_cap_1[4|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[4|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|0] cdac_unit_cap_1[5|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[5|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|0] cdac_unit_cap_1[6|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[6|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|0] cdac_unit_cap_1[7|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[7|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|0] cdac_unit_cap_1[8|0]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[8|0]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|1] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|1] cdac_unit_cap_1[1|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[1|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|1] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|1] cdac_unit_cap_1[3|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[3|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|1] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|1] cdac_unit_cap_1[5|1]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[5|1]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|1] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|1] cdac_unit_cap_1[7|5]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[7|5]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|1] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|2] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|2] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|2] cdac_unit_cap_1[2|6]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|6]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|2] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|2] cdac_unit_cap_1[5|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[5|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|2] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|2] cdac_unit_cap_1[6|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|2] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|2] cdac_unit_cap_1[8|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|3] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|3] cdac_unit_cap_1[1|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[1|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|3] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|3] cdac_unit_cap_1[3|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[3|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|3] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|3] cdac_unit_cap_1[5|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[5|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|3] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|3] cdac_unit_cap_1[7|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[7|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|3] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|4] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|4] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|4] cdac_unit_cap_1[2|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|4] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|4] cdac_unit_cap_1[4|4]/m3_80891_n32882# cdac_unit_cap_1[4|4]/c1_81071_n33152#
+ cdac_unit_cap_1[4|4]/m3_80891_n32882# cdac_unit_cap
Xcdac_unit_cap_1[5|4] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|4] cdac_unit_cap_1[6|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|4] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|4] cdac_unit_cap_1[8|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|5] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|5] cdac_unit_cap_1[1|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[1|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|5] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|5] cdac_unit_cap_1[3|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[3|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|5] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|5] cdac_unit_cap_1[5|5]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[5|5]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|5] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|5] cdac_unit_cap_1[7|5]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[7|5]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|5] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|6] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|6] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|6] cdac_unit_cap_1[2|6]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|6]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|6] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|6] cdac_unit_cap_1[5|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[5|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|6] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|6] cdac_unit_cap_1[6|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|6] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|6] cdac_unit_cap_1[8|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|7] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|7] cdac_unit_cap_1[1|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[1|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|7] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|7] cdac_unit_cap_1[3|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[3|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|7] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|7] cdac_unit_cap_1[5|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[5|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|7] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|7] cdac_unit_cap_1[7|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[7|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|7] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|8] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|8] cdac_unit_cap_1[2|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|8] cdac_unit_cap_1[2|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[2|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|8] cdac_unit_cap_1[4|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|8] cdac_unit_cap_1[4|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[4|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|8] cdac_unit_cap_1[6|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|8] cdac_unit_cap_1[6|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[6|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|8] cdac_unit_cap_1[8|7]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|7]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|8] cdac_unit_cap_1[8|8]/m3_80891_n32882# m4_99908_n7967# cdac_unit_cap_1[8|8]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[0|9] cdac_unit_cap_1[0|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[0|9]/m3_80891_n32882#
+ cdac_unit_cap
Xcdac_unit_cap_1[1|9] cdac_unit_cap_1[1|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[1|9]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[2|9] cdac_unit_cap_1[2|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[2|9]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[3|9] cdac_unit_cap_1[3|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[3|9]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[4|9] cdac_unit_cap_1[4|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[4|9]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[5|9] cdac_unit_cap_1[5|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[5|9]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[6|9] cdac_unit_cap_1[6|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[6|9]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[7|9] cdac_unit_cap_1[7|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[7|9]/c2_81071_n33152#
+ cdac_unit_cap
Xcdac_unit_cap_1[8|9] cdac_unit_cap_1[8|9]/m3_80891_n32882# m4_81638_n9537# cdac_unit_cap_1[8|9]/c2_81071_n33152#
+ cdac_unit_cap
.ends

.subckt cdac_ratioed_cap c1_81071_n33170# m3_80891_n32900# c2_81071_n33170#
X0 c2_81071_n33170# c1_81071_n33170# sky130_fd_pr__cap_mim_m3_2 l=7.055 w=7
X1 c1_81071_n33170# m3_80891_n32900# sky130_fd_pr__cap_mim_m3_1 l=7.055 w=7
.ends

.subckt EF_BANK_CAP_12 D8 D0 D4 VP1 D9 D5 D1 D2 D6 VSS D7 D3 D10 D11 Vref w_58549_n26640#
+ VP2
Xcap_array_half_0 VSS VSS D8 D11 VSS VSS D11 VSS D7 VSS VSS D9 VSS VSS VSS VSS VSS
+ D8 VSS D9 VSS VSS VSS VSS VSS D10 VSS VSS D10 D9 D10 VSS VSS D6 VSS D10 D11 VSS
+ VSS VSS VSS VSS VSS VP2 D7 VSS VSS VSS VSS VP2 VSS VSS VSS D11 cap_array_half
Xcap_array_half_1 VSS VSS D2 D5 VSS VSS D5 VSS D1 VSS VSS D3 VSS VSS VSS Vref VSS
+ D2 VSS D3 VSS VSS VSS VSS VSS D4 VP1 VSS D4 D3 D4 VSS VSS D0 VSS D4 D5 VSS VSS VSS
+ VSS VSS VSS VP1 D1 VSS VSS VSS VSS VP1 VSS VSS VSS D5 cap_array_half
Xcdac_ratioed_cap_0[0] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[1] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[2] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[3] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[4] VP1 VP2 VP2 cdac_ratioed_cap
Xcdac_ratioed_cap_0[5] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[6] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[7] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[8] VSS VSS VSS cdac_ratioed_cap
Xcdac_ratioed_cap_0[9] VSS VSS VSS cdac_ratioed_cap
.ends

.subckt cdac_lvlshift_array HOLD RST SEL0 SEL1 SEL2 SEL3 SEL4 SEL5 SEL6 SEL7 SEL8
+ SEL9 SEL10 SEL11 HOLD_3P3 RST_3P3 SEL0_3P3 SEL1_3P3 SEL2_3P3 SEL3_3P3 SEL5_3P3 SEL6_3P3
+ SEL7_3P3 SEL8_3P3 SEL9_3P3 SEL10_3P3 SEL11_3P3 VDD3P3 VDD1P8 HOLDB_3P3 SEL4_3P3
+ VSS
Xsky130_fd_sc_hvl__decap_4_7 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__decap_4_8 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__decap_4_9 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__inv_2_0 HOLD_3P3 VSS VSS VDD3P3 VDD3P3 HOLDB_3P3 sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_10 SEL8 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 SEL0 VDD1P8 VSS VDD3P3 VDD3P3 SEL0_3P3 VDD3P3 VSS
+ VSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__diode_2_11 SEL10 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_1 HOLD VDD1P8 VSS VDD3P3 VDD3P3 HOLD_3P3 VDD3P3 VSS
+ VSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__diode_2_12 SEL9 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_2 RST VDD1P8 VSS VDD3P3 VDD3P3 RST_3P3 VDD3P3 VSS
+ VSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__diode_2_13 SEL11 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_3 SEL2 VDD1P8 VSS VDD3P3 VDD3P3 SEL2_3P3 VDD3P3 VSS
+ VSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_4 SEL1 VDD1P8 VSS VDD3P3 VDD3P3 SEL1_3P3 VDD3P3 VSS
+ VSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_5 SEL3 VDD1P8 VSS VDD3P3 VDD3P3 SEL3_3P3 VDD3P3 VSS
+ VSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_7 SEL5 VDD1P8 VSS VDD3P3 VDD3P3 SEL5_3P3 VDD3P3 VSS
+ VSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_6 SEL4 VDD1P8 VSS VDD3P3 VDD3P3 SEL4_3P3 VDD3P3 VSS
+ VSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_8 SEL6 VDD1P8 VSS VDD3P3 VDD3P3 SEL6_3P3 VDD3P3 VSS
+ VSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_9 SEL7 VDD1P8 VSS VDD3P3 VDD3P3 SEL7_3P3 VDD3P3 VSS
+ VSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__decap_4_10 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__decap_4_11 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_0 SEL1 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_13 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__decap_4_12 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__lsbuflv2hv_1_10 SEL9 VDD1P8 VSS VDD3P3 VDD3P3 SEL9_3P3 VDD3P3 VSS
+ VSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__diode_2_1 HOLD VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_11 SEL8 VDD1P8 VSS VDD3P3 VDD3P3 SEL8_3P3 VDD3P3 VSS
+ VSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__diode_2_2 RST VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_14 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__lsbuflv2hv_1_12 SEL10 VDD1P8 VSS VDD3P3 VDD3P3 SEL10_3P3 VDD3P3
+ VSS VSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__diode_2_3 SEL0 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_13 SEL11 VDD1P8 VSS VDD3P3 VDD3P3 SEL11_3P3 VDD3P3
+ VSS VSS sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__diode_2_4 SEL2 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_5 SEL3 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_6 SEL4 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_0 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_7 SEL7 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_8 SEL5 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_1 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_9 SEL6 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_2 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__decap_4_3 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__decap_4_5 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__decap_4_4 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__decap_4_6 VSS VSS VDD3P3 VDD3P3 sky130_fd_sc_hvl__decap_4
.ends

.subckt sky130_ef_ip__cdac3v_12bit SELD2 SELD3 SELD4 SELD5 SELD6 SELD7 SELD8 SELD9
+ VDD DVDD OUT RST SELD10 SELD11 OUTNC SELD0 SELD1 Vref VIN HOLD VCM VL VH VSS DVSS
Xx1 OUT OUTNC VDD DVDD VSS x1/HOLD DVSS x1/HOLDB VIN DVDD VSS EF_SW_RST
Xx3 x3/SELD2 x3/SELD3 x3/SELD0 x3/SELD1 x3/SELD4 x4/D1 x3/SELD5 x3/SELD9 x3/SELD8
+ x4/D5 x3/SELD7 x4/D9 x3/SELD6 x4/D8 x4/D7 DVSS x3/SELD10 x3/SELD11 VCM x4/D11 x4/D0
+ cdac_lvlshift_array_0/RST_3P3 x4/D4 x4/D2 cdac_lvlshift_array_0/RST_3P3 x4/D10 VH
+ DVDD x4/D6 x4/D3 VDD VL VSS EF_AMUX0201_ARRAY1
Xx4 x4/D8 x4/D0 x4/D4 OUTNC x4/D9 x4/D5 x4/D1 x4/D2 x4/D6 VSS x4/D7 x4/D3 x4/D10 x4/D11
+ Vref VDD OUT EF_BANK_CAP_12
Xcdac_lvlshift_array_0 HOLD RST SELD0 SELD1 SELD2 SELD3 SELD4 SELD5 SELD6 SELD7 SELD8
+ SELD9 SELD10 SELD11 x1/HOLD cdac_lvlshift_array_0/RST_3P3 x3/SELD0 x3/SELD1 x3/SELD2
+ x3/SELD3 x3/SELD5 x3/SELD6 x3/SELD7 x3/SELD8 x3/SELD9 x3/SELD10 x3/SELD11 VDD DVDD
+ x1/HOLDB x3/SELD4 DVSS cdac_lvlshift_array
.ends

.subckt sky130_fd_pr__res_high_po_0p35_AW5QUD a_n35_300# a_n35_n732# VSUBS
X0 a_n35_300# a_n35_n732# VSUBS sky130_fd_pr__res_high_po_0p35 l=3.16
.ends

.subckt dac_3v_cell m1_814_1199# w_318_n275# m1_545_847# m1_387_847# m1_824_799# m1_290_1114#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS m1_545_212# m1_663_847# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732#
+ m1_300_n125# m1_821_212# m1_814_483# m1_663_212# m1_814_591# w_316_892# m1_814_n125#
+ m1_290_591# sky130_fd_pr__res_high_po_0p35_AW5QUD_0/a_n35_300# m1_155_n223# m1_290_344#
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_0 sky130_fd_pr__res_high_po_0p35_AW5QUD_0/a_n35_300#
+ m1_155_n223# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_1 m1_824_799# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_545_847# m1_387_847# m1_290_1114# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_663_847# m1_814_1199# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_821_212# m1_663_212# m1_814_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# m1_300_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# m1_290_591# m1_545_847# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_663_847# m1_814_591# m1_824_799# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# m1_290_344# m1_545_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_663_212# m1_814_483# m1_821_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
.ends

.subckt dac_3v_cell_top m1_814_1199# w_318_n275# m1_545_847# m1_387_847# m1_824_799#
+ w_318_892# m1_290_1114# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS m1_545_212#
+ m1_663_847# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732# m1_300_n125# m4_97_801#
+ m1_821_212# m4_97_1059# m1_814_483# m1_663_212# m1_814_591# m1_814_n125# m1_290_591#
+ m1_155_n223# m1_290_344#
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_0 m1_824_799# m1_155_n223# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_1 m1_824_799# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_545_847# m1_387_847# m1_290_1114# w_318_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_663_847# m1_814_1199# w_318_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_821_212# m1_663_212# m1_814_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# m1_300_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# m1_290_591# m1_545_847# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_663_847# m1_814_591# m1_824_799# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# m1_290_344# m1_545_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_663_212# m1_814_483# m1_821_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
.ends

.subckt dac_3v_cell_odd m1_814_1199# w_318_n275# m1_545_847# m1_387_847# m1_824_799#
+ m1_290_1114# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS m1_545_212# m1_663_847#
+ m1_155_n223# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732# m1_300_n125# m1_821_212#
+ m1_814_483# m1_663_212# m1_814_591# w_316_892# m1_814_n125# m1_290_591# sky130_fd_pr__res_high_po_0p35_AW5QUD_0/a_n35_300#
+ m1_290_344#
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_0 sky130_fd_pr__res_high_po_0p35_AW5QUD_0/a_n35_300#
+ m1_155_n223# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_1 m1_824_799# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_545_847# m1_387_847# m1_290_1114# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_663_847# m1_814_1199# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_821_212# m1_663_212# m1_814_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# m1_300_n125# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# m1_290_591# m1_545_847# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_663_847# m1_814_591# m1_824_799# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# m1_290_344# m1_545_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_663_212# m1_814_483# m1_821_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
.ends

.subckt dac_3v_column_odd m3_31_13582# res_in0 b3_uq0 b0_uq0 b0_uq5 dac_3v_cell_top_0/m4_97_801#
+ b0_uq4 b0_uq11 b2b_uq0 b4 b4b b0b_uq13 b2 b0_uq10 b1_uq5 dac_3v_cell_0[2]/w_316_892#
+ dac_3v_cell_0[1]/w_316_892# b1_uq4 b0 dac_3v_cell_top_0/m4_97_1059# b1_uq6 b0_uq12
+ b0b_uq6 b0b_uq5 m3_30_13212# b0b_uq4 b1_uq0 b0b_uq3 b3b_uq0 b2b_uq2 b0b_uq2 b0b_uq1
+ b0_uq14 b0b_uq14 dac_3v_cell_0[0]/w_316_892# b0b_uq11 b0b_uq0 b0_uq1 b0_uq6 b0b_uq10
+ out_5 b1_uq1 b1 b3b m2_791_14877# m2_801_196# dum_in0 b0b_uq12 b1b_uq6 res_out1
+ b0_uq13 b2_uq2 b2b_uq1 out4 b1b_uq5 dac_3v_cell_0[4]/w_316_892# b2_uq1 b3 dac_3v_cell_odd_0/w_316_892#
+ b1b_uq4 b0_uq3 b2_uq0 b1b_uq3 b1b_uq2 b1b_uq1 b0_uq2 b1_uq2 b1b_uq0 b0b_uq9 m2_791_1314#
+ dac_3v_cell_0[5]/w_316_892# b0_uq9 in_5 b0b dum_out1 b1_uq3 b0_uq8 dac_3v_cell_0[3]/w_316_892#
+ b1b b0b_uq8 b0b_uq7 b0_uq7 m2_801_13759# b2b VSUBS
Xdac_3v_cell_0[0] b0_uq2 dac_3v_cell_odd_0/w_316_892# out0_2 out0_1_0 dac_3v_cell_0[0]/m1_824_799#
+ b2b_uq0 VSUBS out0_0_0 out1_0_3 dac_3v_cell_odd_0/m1_824_799# b0b_uq1 out1_1_1 b1b
+ out1_0_3 b0b_uq2 dac_3v_cell_0[0]/w_316_892# b1 b2_uq0 dac_3v_cell_0[1]/m1_155_n223#
+ dac_3v_cell_0[0]/m1_155_n223# b0_uq1 dac_3v_cell
Xdac_3v_cell_0[1] b0b_uq4 dac_3v_cell_0[0]/w_316_892# out0_0_1 out0_1_0 dac_3v_cell_0[1]/m1_824_799#
+ b1_uq1 VSUBS out0_0_1 out1_0_2 dac_3v_cell_0[0]/m1_824_799# b0_uq3 out1_1_1 b2b
+ out1_2 b0_uq4 dac_3v_cell_0[1]/w_316_892# b2 b1b_uq1 dac_3v_cell_0[2]/m1_155_n223#
+ dac_3v_cell_0[1]/m1_155_n223# b0b_uq3 dac_3v_cell
Xdac_3v_cell_0[2] b0_uq6 dac_3v_cell_0[1]/w_316_892# out_3 out0_2 dac_3v_cell_0[2]/m1_824_799#
+ b3b_uq0 VSUBS out0_0_1 out1_0_2 dac_3v_cell_0[1]/m1_824_799# b0b_uq5 out1_1_1 b1_uq2
+ out1_0_2 b0b_uq6 dac_3v_cell_0[2]/w_316_892# b1b_uq2 b3_uq0 dac_3v_cell_0[3]/m1_155_n223#
+ dac_3v_cell_0[2]/m1_155_n223# b0_uq5 dac_3v_cell
Xdac_3v_cell_0[3] b0b_uq8 dac_3v_cell_0[2]/w_316_892# out0_0_2 m3_296_8710# dac_3v_cell_0[3]/m1_824_799#
+ b1b_uq3 VSUBS out0_0_2 out1_0_1 dac_3v_cell_0[2]/m1_824_799# b0_uq7 out1_2 b3b out_3
+ b0_uq8 dac_3v_cell_0[3]/w_316_892# b3 b1_uq3 dac_3v_cell_0[4]/m1_155_n223# dac_3v_cell_0[3]/m1_155_n223#
+ b0b_uq7 dac_3v_cell
Xdac_3v_cell_0[4] b0_uq10 dac_3v_cell_0[3]/w_316_892# out0_2 m3_296_8710# dac_3v_cell_0[4]/m1_824_799#
+ b2_uq1 VSUBS out0_0_2 out1_0_1 dac_3v_cell_0[3]/m1_824_799# b0b_uq9 out1_1_0 b1b_uq4
+ out1_0_1 b0b_uq10 dac_3v_cell_0[4]/w_316_892# b1_uq4 b2b_uq1 dac_3v_cell_0[5]/m1_155_n223#
+ dac_3v_cell_0[4]/m1_155_n223# b0_uq9 dac_3v_cell
Xdac_3v_cell_0[5] b0b_uq12 dac_3v_cell_0[4]/w_316_892# out0_0_3 m3_296_8710# dac_3v_cell_0[5]/m1_824_799#
+ b1_uq5 VSUBS out0_0_3 out1_0_0 dac_3v_cell_0[4]/m1_824_799# b0_uq11 out1_1_0 b2_uq2
+ out1_2 b0_uq12 dac_3v_cell_0[5]/w_316_892# b2b_uq2 b1b_uq5 dac_3v_cell_top_0/m1_155_n223#
+ dac_3v_cell_0[5]/m1_155_n223# b0b_uq11 dac_3v_cell
Xdac_3v_cell_1 m2_791_1314# m2_801_196# m2_329_1119# m2_329_1119# res_out1 m2_791_1314#
+ VSUBS m2_457_485# m2_329_1119# dum_out1 m2_801_196# m2_457_485# VSUBS m2_457_485#
+ VSUBS m2_791_1314# m2_801_196# VSUBS res_in0 dum_in0 VSUBS dac_3v_cell
Xdac_3v_cell_2 m2_791_14877# m2_801_13759# m2_331_14682# m2_331_14682# dum_out0 m2_791_14877#
+ VSUBS m2_458_14048# m2_331_14682# res_in1 m2_801_13759# m2_458_14048# VSUBS m2_458_14048#
+ VSUBS m2_791_14877# m2_801_13759# VSUBS dum_out0 res_in1 VSUBS dac_3v_cell
Xdac_3v_cell_top_0 b0_uq14 dac_3v_cell_0[5]/w_316_892# in_5 out_5 res_in1 m2_801_13759#
+ m3_31_13582# VSUBS out0_0_3 out1_0_0 dac_3v_cell_0[5]/m1_824_799# b0b_uq13 dac_3v_cell_top_0/m4_97_801#
+ out1_1_0 dac_3v_cell_top_0/m4_97_1059# b1_uq6 out1_0_0 b0b_uq14 b1b_uq6 m3_30_13212#
+ dac_3v_cell_top_0/m1_155_n223# b0_uq13 dac_3v_cell_top
Xdac_3v_cell_odd_0 b0b m2_791_1314# out0_0_0 out0_1_0 dac_3v_cell_odd_0/m1_824_799#
+ b1b_uq0 VSUBS out0_0_0 out1_0_3 res_in0 res_out1 b0_uq0 out_3 b4 out4 b0 dac_3v_cell_odd_0/w_316_892#
+ b4b b1_uq0 dac_3v_cell_0[0]/m1_155_n223# b0b_uq0 dac_3v_cell_odd
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AQ2WAW a_1293_n197# a_n761_n197# a_1235_n100#
+ a_n1551_n197# a_761_n100# a_n29_n100# a_1393_n100# a_1451_n197# a_n187_n100# a_1551_n100#
+ a_n819_n100# a_n345_n100# a_n1609_n100# a_29_n197# a_n977_n100# a_n1135_n100# a_n129_n197#
+ a_187_n197# a_129_n100# a_n503_n100# a_n1293_n100# a_n287_n197# a_819_n197# a_n661_n100#
+ a_345_n197# a_n1077_n197# a_287_n100# a_n1451_n100# a_n919_n197# a_977_n197# a_n445_n197#
+ a_919_n100# a_503_n197# a_n1235_n197# a_445_n100# w_n1809_n397# a_1077_n100# a_1135_n197#
+ a_n603_n197# a_n1393_n197# a_661_n197# a_603_n100#
X0 a_919_n100# a_819_n197# a_761_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_445_n100# a_345_n197# a_287_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_603_n100# a_503_n197# a_445_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_n1293_n100# a_n1393_n197# a_n1451_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_n1451_n100# a_n1551_n197# a_n1609_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X5 a_n977_n100# a_n1077_n197# a_n1135_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_n1135_n100# a_n1235_n197# a_n1293_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 a_n661_n100# a_n761_n197# a_n819_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 a_129_n100# a_29_n197# a_n29_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X9 a_n187_n100# a_n287_n197# a_n345_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X10 a_n819_n100# a_n919_n197# a_n977_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 a_n345_n100# a_n445_n197# a_n503_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X12 a_n503_n100# a_n603_n197# a_n661_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X13 a_n29_n100# a_n129_n197# a_n187_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X14 a_1393_n100# a_1293_n197# a_1235_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X15 a_1077_n100# a_977_n197# a_919_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X16 a_1551_n100# a_1451_n197# a_1393_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X17 a_761_n100# a_661_n197# a_603_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X18 a_287_n100# a_187_n197# a_129_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X19 a_1235_n100# a_1135_n197# a_1077_n100# w_n1809_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UNEQFS a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLJMY6 a_n208_n197# a_208_n100# a_n50_n197# a_50_n100#
+ a_n108_n100# w_n466_n397# a_n266_n100# a_108_n197#
X0 a_208_n100# a_108_n197# a_50_n100# w_n466_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_50_n100# a_n50_n197# a_n108_n100# w_n466_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n108_n100# a_n208_n197# a_n266_n100# w_n466_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_KLWMS5 a_n29_n100# a_n187_n100# w_n545_n397#
+ a_n345_n100# a_29_n197# a_n129_n197# a_187_n197# a_129_n100# a_n287_n197# a_287_n100#
X0 a_129_n100# a_29_n197# a_n29_n100# w_n545_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n187_n100# a_n287_n197# a_n345_n100# w_n545_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X2 a_n29_n100# a_n129_n197# a_n187_n100# w_n545_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_287_n100# a_187_n197# a_129_n100# w_n545_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_HLA228 a_131_1150# a_131_n1582# a_n201_n1582#
+ a_n35_n1582# a_n201_1150# a_n35_1150# a_n331_n1712#
X0 a_n35_1150# a_n35_n1582# a_n331_n1712# sky130_fd_pr__res_xhigh_po_0p35 l=11.66
X1 a_n201_1150# a_n201_n1582# a_n331_n1712# sky130_fd_pr__res_xhigh_po_0p35 l=11.66
X2 a_131_1150# a_131_n1582# a_n331_n1712# sky130_fd_pr__res_xhigh_po_0p35 l=11.66
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_FJGQFC a_n321_n322# a_n29_n100# a_n187_n100#
+ a_129_n100# a_29_n188# a_n129_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n188# a_n187_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_XJGQ2Y a_n321_n322# a_n29_n100# a_n187_n100#
+ a_129_n100# a_29_n188# a_n129_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n29_n100# a_n129_n188# a_n187_n100# a_n321_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_05v0_nvt_BH6ZTK a_n29_n100# a_209_n100# a_n209_n188# a_n401_n322#
+ a_n267_n100# a_29_n188#
X0 a_209_n100# a_29_n188# a_n29_n100# a_n401_n322# sky130_fd_pr__nfet_05v0_nvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.9
X1 a_n29_n100# a_n209_n188# a_n267_n100# a_n401_n322# sky130_fd_pr__nfet_05v0_nvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.9
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Z8JNCQ a_n345_118# a_1393_n2934# a_977_n851#
+ a_603_n1626# a_n1451_2734# a_1551_n2498# a_29_n415# a_n661_554# a_n1551_21# a_1451_1329#
+ a_445_118# a_n445_n851# a_n129_n2595# a_761_554# a_n129_1765# a_n661_2298# a_n187_n754#
+ a_29_n1287# a_n977_n2062# a_345_893# a_287_2298# a_1235_n1626# a_n129_n415# a_977_n3031#
+ a_n1235_n2595# a_445_1862# a_761_n2498# a_n29_n2498# a_603_n318# a_187_1765# a_n503_1426#
+ a_29_2637# a_n1235_n851# a_129_1426# a_919_2734# a_1077_990# a_n287_457# a_187_n415#
+ a_n603_n2595# a_445_n1626# a_n977_990# a_n1293_1426# a_n603_2201# a_1393_n2498#
+ a_n1451_2298# a_1135_2201# a_977_21# a_503_n851# a_919_n1626# a_n1393_2201# a_n1135_n2934#
+ a_n129_2637# a_29_n2159# a_1077_n1626# a_n1609_n2934# a_661_2201# a_187_21# a_n1077_n2595#
+ a_445_2734# a_n187_118# a_1551_n754# a_n503_n2934# a_29_457# a_187_2637# a_129_990#
+ a_287_118# a_1077_1862# a_503_n2595# a_n819_n754# a_n287_1765# a_n445_n2595# a_287_n1626#
+ a_919_2298# a_1235_n318# a_187_893# a_1451_457# a_n287_n415# a_n919_n2595# a_1551_n1626#
+ a_1135_n2595# a_n1551_n2595# a_1451_21# a_n129_n1723# a_n1135_n2498# a_819_1765#
+ a_n603_n851# a_761_n318# a_1135_n851# a_n661_1426# a_n345_n754# a_n1609_n2498# a_819_n415#
+ a_n1393_n851# a_287_1426# a_445_2298# a_n761_2201# a_n919_457# a_n345_n2934# a_n1077_1765#
+ a_n1609_n754# a_n1235_n1723# a_n503_n2498# a_n1609_990# a_1293_2201# a_761_n1626#
+ a_603_1862# a_1077_2734# a_661_n851# a_n29_n1626# a_345_n2595# a_n1235_893# a_n445_21#
+ a_n819_n2934# a_n1077_n415# a_503_457# a_n287_n2595# a_n287_2637# a_345_1765# a_n1451_n2934#
+ a_819_n2595# a_n603_n1723# a_345_n415# a_1393_n1626# a_n1451_1426# a_n1393_n2595#
+ a_n1135_n754# a_819_2637# a_n819_118# a_n129_n1287# a_n29_n318# a_n1551_2201# a_n29_990#
+ a_1235_554# a_n919_1765# a_n1135_554# a_919_118# a_n977_n754# a_1551_990# a_n761_457#
+ a_n187_n2934# a_1393_n318# a_n1077_n1723# a_n1451_990# a_n1077_2637# a_n345_n2498#
+ a_n761_n2595# a_n919_n415# a_1293_457# a_n1235_n1287# a_819_893# a_603_2734# a_187_n2595#
+ a_1077_2298# a_n819_n2498# a_345_2637# a_977_1765# a_n761_n851# a_503_n1723# a_n1293_n2934#
+ a_1235_1862# a_1451_n2595# a_1293_n851# a_n445_n1723# a_n1451_n2498# a_29_1329#
+ a_n1077_21# a_129_n1190# a_n445_1765# a_n603_n1287# a_919_1426# a_977_n415# a_n503_990#
+ a_n919_n1723# a_n661_118# a_n445_n415# a_n129_n2159# a_n661_n2934# a_1135_n1723#
+ a_761_1862# a_603_990# a_n1551_n1723# a_n1135_n1626# a_n129_1329# a_761_118# a_n919_2637#
+ a_n187_n318# a_n1077_893# a_345_457# a_661_n2595# a_n1609_n1626# a_n187_n2498# a_345_21#
+ a_n1077_n1287# a_661_893# a_29_21# a_n503_n754# a_n1235_n2159# a_n1551_n851# a_445_1426#
+ a_603_2298# a_129_n754# a_n503_n1626# a_n1235_1765# a_603_n1190# a_n1293_n754# a_187_1329#
+ a_1451_2201# a_977_2637# a_345_n1723# a_1293_n2595# a_1235_2734# a_n287_n1723# a_n1293_n2498#
+ a_503_n1287# a_n1235_n415# a_129_n2062# a_n445_n1287# a_n129_893# a_n445_2637# a_n977_554#
+ a_1077_554# a_n603_n2159# a_503_1765# a_819_n1723# a_1393_990# a_1235_n1190# a_n1293_990#
+ a_n919_n1287# a_503_n415# a_n29_1862# a_761_2734# a_n1393_n1723# a_1135_n1287# a_n661_n2498#
+ a_n1551_n1287# a_n977_n2934# a_1393_1862# a_n1077_n2159# a_977_n2595# a_n761_n1723#
+ a_1551_n318# a_n345_n1626# a_445_n1190# a_603_n2062# a_n1235_2637# a_n345_990# a_129_554#
+ a_187_n1723# a_1077_1426# a_345_n1287# a_n603_21# a_n819_n1626# a_503_n2159# a_919_n1190#
+ a_1235_2298# a_445_990# a_n819_n318# a_n287_n1287# a_n287_1329# a_n445_n2159# a_29_n3031#
+ a_503_2637# a_1451_n1723# a_n1451_n1626# a_187_457# a_819_n1287# a_1451_n851# a_1077_n1190#
+ a_1235_n2062# a_n919_n2159# a_n603_1765# a_n661_n754# a_1135_1765# a_n29_2734# a_n1393_n1287#
+ a_1135_n2159# a_761_2298# a_287_n754# a_n1551_n2159# a_819_1329# a_n187_1862# a_n1393_1765#
+ a_n603_n415# a_1135_n415# a_1393_2734# a_n977_n2498# a_n1393_n415# a_n345_n318#
+ a_661_n1723# a_661_1765# a_n187_n1626# a_n1609_n318# a_287_n1190# a_445_n2062# a_n1077_1329#
+ a_n761_n1287# a_n1609_554# a_603_1426# a_187_n1287# a_n1235_457# a_661_n415# a_345_n2159#
+ a_1551_n1190# a_919_n2062# a_n287_n2159# a_n1451_n754# a_345_1329# a_1293_n1723#
+ a_n1551_893# a_n1293_n1626# a_1451_n1287# a_819_n2159# a_1077_n2062# a_n603_2637#
+ a_n1235_21# a_1135_2637# a_n29_2298# a_n1135_n318# a_n1393_n2159# a_n187_2734# a_n1393_2637#
+ a_n187_990# a_n661_n1626# a_761_n1190# a_n29_554# a_1235_118# a_n919_1329# a_1393_2298#
+ a_n1135_118# a_n977_n318# a_n29_n1190# a_287_990# a_661_n1287# a_n603_893# a_661_2637#
+ a_1551_554# a_287_n2062# a_n1451_554# a_1551_1862# a_n761_n2159# a_1135_893# a_503_21#
+ a_977_n1723# a_819_457# a_n761_1765# a_187_n2159# a_1293_1765# a_1393_n1190# a_1551_n2062#
+ a_919_n754# a_n819_1862# a_n761_n415# a_977_1329# a_1293_n1287# a_1235_1426# a_1451_n2159#
+ a_1293_n415# a_n445_1329# a_n503_554# a_n187_2298# a_761_1426# a_603_554# a_761_n2062#
+ a_n1077_457# a_445_n754# a_n29_n2062# a_n345_1862# a_n1551_1765# a_n977_n1626# a_661_n2159#
+ a_n1393_893# a_1551_2734# a_n1609_1862# a_29_2201# a_661_457# a_n1551_n415# a_n503_n318#
+ a_n761_2637# a_977_n1287# a_129_n318# a_1393_n2062# a_1293_2637# a_n1235_1329# a_n819_2734#
+ a_n1293_n318# a_n129_n3031# a_1293_n2159# a_n129_457# a_n129_2201# a_1077_118# a_n819_990#
+ a_n977_118# a_n1135_n1190# a_503_1329# a_n445_893# a_1393_554# a_919_990# a_n1135_1862#
+ a_n1293_554# a_1135_21# a_n1609_n1190# a_n1235_n3031# a_n29_1426# a_n919_21# a_n345_2734#
+ a_n1551_2637# a_n503_n1190# a_977_893# a_n977_1862# a_187_2201# a_1393_1426# a_n1609_2734#
+ a_1551_2298# a_1077_n754# a_n761_21# a_977_n2159# a_n603_n3031# a_n129_21# a_n345_554#
+ a_129_118# a_n819_2298# a_29_n851# a_1451_1765# a_n661_990# a_445_554# a_n1135_n2062#
+ a_129_n2934# a_761_990# a_1451_n415# a_n1135_2734# a_n1077_n3031# a_n603_1329# a_n661_n318#
+ a_n1609_n2062# a_1135_1329# a_n129_n851# a_287_n318# a_n187_1426# a_n1393_1329#
+ a_n345_n1190# a_n503_n2062# a_n977_2734# a_n345_2298# a_503_n3031# a_603_n754# a_n1609_2298#
+ a_n287_2201# a_n819_n1190# a_n445_n3031# a_n503_1862# a_661_1329# a_129_1862# a_n1609_118#
+ a_n1451_n1190# a_187_n851# a_n287_893# a_603_n2934# a_n1293_1862# a_n919_n3031#
+ a_n1393_21# a_1451_2637# a_1135_n3031# a_n1551_n3031# a_n1451_n318# a_819_2201#
+ a_n1551_457# a_129_n2498# a_29_n2595# a_n1135_2298# a_1235_n2934# a_819_21# a_n1077_2201#
+ a_n187_n1190# a_n345_n2062# a_n187_554# a_n977_2298# a_661_21# w_n1809_n3231# a_n29_118#
+ a_345_n3031# a_29_893# a_n819_n2062# a_n287_n3031# a_n503_2734# a_n603_457# a_287_554#
+ a_345_2201# a_1551_118# a_n1451_118# a_1551_1426# a_129_2734# a_n1293_n1190# a_819_n3031#
+ a_1135_457# a_n1451_n2062# a_445_n2934# a_n1293_2734# a_1235_n754# a_n761_1329#
+ a_603_n2498# a_1451_893# a_1293_1329# a_919_n318# a_n287_n851# a_n1393_n3031# a_n819_1426#
+ a_919_n2934# a_n661_n1190# a_n919_2201# a_761_n754# a_1077_n2934# a_n661_1862# a_1235_n2498#
+ a_n503_118# a_819_n851# a_287_1862# a_n761_n3031# a_n187_n2062# a_603_118# a_187_n3031#
+ a_n919_893# a_445_n318# a_n345_1426# a_n1551_1329# a_n503_2298# a_977_2201# a_n1393_457#
+ a_n1077_n851# a_1451_n3031# a_503_893# a_n1609_1426# a_n1293_n2062# a_287_n2934#
+ a_129_2298# a_n445_2201# a_445_n2498# a_n1293_2298# a_345_n851# a_1551_n2934# a_n1451_1862#
+ a_919_n2498# a_1293_21# a_n819_554# a_n661_n2062# a_n29_n754# a_129_n1626# a_n661_2734#
+ a_29_n1723# a_661_n3031# a_1077_n2498# a_1235_990# a_n445_457# a_919_554# a_1393_118#
+ a_n1135_990# a_n977_n1190# a_n1135_1426# a_287_2734# a_n1293_118# a_n761_893# a_1393_n754#
+ a_n919_n851# a_761_n2934# a_1293_893# a_n1235_2201# a_977_457# a_n977_1426# a_n29_n2934#
+ a_n287_21# a_1293_n3031# a_1077_n318# a_287_n2498# a_503_2201# a_29_1765# a_919_1862#
X0 a_919_n2934# a_819_n3031# a_761_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_1077_n1626# a_977_n1723# a_919_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 a_n1451_n1626# a_n1551_n1723# a_n1609_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 a_919_n1190# a_819_n1287# a_761_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 a_287_554# a_187_457# a_129_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 a_1393_990# a_1293_893# a_1235_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X6 a_n29_n754# a_n129_n851# a_n187_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 a_603_n754# a_503_n851# a_445_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 a_129_n2062# a_29_n2159# a_n29_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X9 a_1235_1862# a_1135_1765# a_1077_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X10 a_1235_554# a_1135_457# a_1077_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 a_n1135_1862# a_n1235_1765# a_n1293_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X12 a_1077_n2934# a_977_n3031# a_919_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X13 a_n1451_n2934# a_n1551_n3031# a_n1609_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X14 a_1077_990# a_977_893# a_919_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X15 a_n1451_n1190# a_n1551_n1287# a_n1609_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X16 a_919_n2498# a_819_n2595# a_761_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X17 a_1077_n1190# a_977_n1287# a_919_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X18 a_n345_n1626# a_n445_n1723# a_n503_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X19 a_919_554# a_819_457# a_761_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X20 a_1551_990# a_1451_893# a_1393_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X21 a_445_554# a_345_457# a_287_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X22 a_n1293_118# a_n1393_21# a_n1451_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X23 a_445_n2062# a_345_n2159# a_287_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X24 a_n819_1426# a_n919_1329# a_n977_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X25 a_1077_n2498# a_977_n2595# a_919_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X26 a_n1451_n2498# a_n1551_n2595# a_n1609_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X27 a_n345_n2934# a_n445_n3031# a_n503_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X28 a_n345_n1190# a_n445_n1287# a_n503_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X29 a_n1135_n754# a_n1235_n851# a_n1293_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X30 a_1235_n754# a_1135_n851# a_1077_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X31 a_n661_1426# a_n761_1329# a_n819_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X32 a_761_990# a_661_893# a_603_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X33 a_n819_n1626# a_n919_n1723# a_n977_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X34 a_603_554# a_503_457# a_445_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X35 a_n819_2734# a_n919_2637# a_n977_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X36 a_n1451_118# a_n1551_21# a_n1609_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X37 a_n977_n1626# a_n1077_n1723# a_n1135_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X38 a_919_n2062# a_819_n2159# a_761_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X39 a_919_1426# a_819_1329# a_761_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X40 a_n345_n2498# a_n445_n2595# a_n503_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X41 a_1235_n1626# a_1135_n1723# a_1077_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X42 a_n661_2734# a_n761_2637# a_n819_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X43 a_287_990# a_187_893# a_129_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X44 a_n819_n2934# a_n919_n3031# a_n977_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X45 a_n819_n318# a_n919_n415# a_n977_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X46 a_n819_n1190# a_n919_n1287# a_n977_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X47 a_1235_990# a_1135_893# a_1077_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X48 a_n977_118# a_n1077_21# a_n1135_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X49 a_n819_2298# a_n919_2201# a_n977_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X50 a_n187_1426# a_n287_1329# a_n345_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X51 a_761_1426# a_661_1329# a_603_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X52 a_n977_n2934# a_n1077_n3031# a_n1135_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X53 a_1077_n2062# a_977_n2159# a_919_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X54 a_n977_n1190# a_n1077_n1287# a_n1135_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X55 a_n1451_n2062# a_n1551_n2159# a_n1609_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X56 a_919_2734# a_819_2637# a_761_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X57 a_n661_n318# a_n761_n415# a_n819_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X58 a_1235_n2934# a_1135_n3031# a_1077_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X59 a_1393_n1626# a_1293_n1723# a_1235_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X60 a_n661_2298# a_n761_2201# a_n819_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X61 a_919_990# a_819_893# a_761_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X62 a_n819_n2498# a_n919_n2595# a_n977_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X63 a_603_n1626# a_503_n1723# a_445_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X64 a_1235_n1190# a_1135_n1287# a_1077_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X65 a_445_990# a_345_893# a_287_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X66 a_n1293_554# a_n1393_457# a_n1451_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X67 a_n187_2734# a_n287_2637# a_n345_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X68 a_761_2734# a_661_2637# a_603_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X69 a_n819_1862# a_n919_1765# a_n977_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X70 a_n1135_118# a_n1235_21# a_n1293_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X71 a_919_n318# a_819_n415# a_761_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X72 a_n977_n2498# a_n1077_n2595# a_n1135_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X73 a_1393_n2934# a_1293_n3031# a_1235_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X74 a_919_2298# a_819_2201# a_761_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X75 a_n345_n2062# a_n445_n2159# a_n503_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X76 a_1393_n1190# a_1293_n1287# a_1235_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X77 a_287_1426# a_187_1329# a_129_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X78 a_603_n2934# a_503_n3031# a_445_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X79 a_1235_n2498# a_1135_n2595# a_1077_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X80 a_761_n1626# a_661_n1723# a_603_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X81 a_603_n1190# a_503_n1287# a_445_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X82 a_n661_1862# a_n761_1765# a_n819_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X83 a_n187_n318# a_n287_n415# a_n345_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X84 a_761_n318# a_661_n415# a_603_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X85 a_n1293_1426# a_n1393_1329# a_n1451_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X86 a_1393_1426# a_1293_1329# a_1235_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X87 a_603_990# a_503_893# a_445_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X88 a_n187_2298# a_n287_2201# a_n345_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X89 a_761_2298# a_661_2201# a_603_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X90 a_n1451_554# a_n1551_457# a_n1609_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X91 a_287_2734# a_187_2637# a_129_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X92 a_761_n2934# a_661_n3031# a_603_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X93 a_1393_n2498# a_1293_n2595# a_1235_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X94 a_919_1862# a_819_1765# a_761_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X95 a_761_n1190# a_661_n1287# a_603_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X96 a_n661_118# a_n761_21# a_n819_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X97 a_603_n2498# a_503_n2595# a_445_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X98 a_n819_n2062# a_n919_n2159# a_n977_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X99 a_1393_2734# a_1293_2637# a_1235_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X100 a_n1293_2734# a_n1393_2637# a_n1451_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X101 a_n819_n754# a_n919_n851# a_n977_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X102 a_n977_554# a_n1077_457# a_n1135_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X103 a_129_118# a_29_21# a_n29_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X104 a_n187_1862# a_n287_1765# a_n345_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X105 a_761_1862# a_661_1765# a_603_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X106 a_287_n318# a_187_n415# a_129_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X107 a_n977_n2062# a_n1077_n2159# a_n1135_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X108 a_287_2298# a_187_2201# a_129_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X109 a_n661_n754# a_n761_n851# a_n819_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X110 a_761_n2498# a_661_n2595# a_603_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X111 a_n187_118# a_n287_21# a_n345_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X112 a_1393_n318# a_1293_n415# a_1235_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X113 a_1235_n2062# a_1135_n2159# a_1077_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X114 a_n1293_n318# a_n1393_n415# a_n1451_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X115 a_1393_2298# a_1293_2201# a_1235_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X116 a_n1293_2298# a_n1393_2201# a_n1451_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X117 a_n345_1426# a_n445_1329# a_n503_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X118 a_n1293_990# a_n1393_893# a_n1451_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X119 a_n503_n1626# a_n603_n1723# a_n661_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X120 a_n1135_554# a_n1235_457# a_n1293_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X121 a_919_n754# a_819_n851# a_761_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X122 a_1393_n2062# a_1293_n2159# a_1235_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X123 a_n819_118# a_n919_21# a_n977_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X124 a_287_n1626# a_187_n1723# a_129_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X125 a_287_1862# a_187_1765# a_129_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X126 a_603_n2062# a_503_n2159# a_445_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X127 a_n345_2734# a_n445_2637# a_n503_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X128 a_129_1426# a_29_1329# a_n29_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X129 a_n345_118# a_n445_21# a_n503_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X130 a_n187_n754# a_n287_n851# a_n345_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X131 a_761_n754# a_661_n851# a_603_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X132 a_n661_n1626# a_n761_n1723# a_n819_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X133 a_n1293_1862# a_n1393_1765# a_n1451_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X134 a_1393_1862# a_1293_1765# a_1235_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X135 a_n503_n2934# a_n603_n3031# a_n661_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X136 a_n1451_990# a_n1551_893# a_n1609_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X137 a_n503_n1190# a_n603_n1287# a_n661_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X138 a_445_1426# a_345_1329# a_287_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X139 a_287_n2934# a_187_n3031# a_129_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X140 a_761_n2062# a_661_n2159# a_603_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X141 a_n345_n318# a_n445_n415# a_n503_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X142 a_287_n1190# a_187_n1287# a_129_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X143 a_129_2734# a_29_2637# a_n29_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X144 a_1551_1426# a_1451_1329# a_1393_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X145 a_n661_554# a_n761_457# a_n819_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X146 a_n345_2298# a_n445_2201# a_n503_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X147 a_n1451_1426# a_n1551_1329# a_n1609_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X148 a_n661_n2934# a_n761_n3031# a_n819_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X149 a_n1135_n1626# a_n1235_n1723# a_n1293_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X150 a_n503_118# a_n603_21# a_n661_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X151 a_n503_n2498# a_n603_n2595# a_n661_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X152 a_n661_n1190# a_n761_n1287# a_n819_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X153 a_n977_990# a_n1077_893# a_n1135_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X154 a_129_554# a_29_457# a_n29_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X155 a_445_2734# a_345_2637# a_287_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X156 a_287_n754# a_187_n851# a_129_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X157 a_129_n318# a_29_n415# a_n29_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X158 a_287_n2498# a_187_n2595# a_129_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X159 a_n1451_2734# a_n1551_2637# a_n1609_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X160 a_1551_2734# a_1451_2637# a_1393_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X161 a_129_2298# a_29_2201# a_n29_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X162 a_n187_554# a_n287_457# a_n345_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X163 a_1393_n754# a_1293_n851# a_1235_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X164 a_n1293_n754# a_n1393_n851# a_n1451_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X165 a_n1135_n2934# a_n1235_n3031# a_n1293_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X166 a_n1293_n1626# a_n1393_n1723# a_n1451_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X167 a_n29_118# a_n129_21# a_n187_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X168 a_445_n318# a_345_n415# a_287_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X169 a_n1135_n1190# a_n1235_n1287# a_n1293_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X170 a_n661_n2498# a_n761_n2595# a_n819_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X171 a_n345_1862# a_n445_1765# a_n503_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X172 a_1551_n1626# a_1451_n1723# a_1393_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X173 a_n29_n1626# a_n129_n1723# a_n187_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X174 a_445_2298# a_345_2201# a_287_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X175 a_n977_1426# a_n1077_1329# a_n1135_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X176 a_n1135_990# a_n1235_893# a_n1293_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X177 a_n1451_n318# a_n1551_n415# a_n1609_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X178 a_1551_n318# a_1451_n415# a_1393_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X179 a_1077_1426# a_977_1329# a_919_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X180 a_n819_554# a_n919_457# a_n977_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X181 a_1393_118# a_1293_21# a_1235_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X182 a_n1293_n2934# a_n1393_n3031# a_n1451_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X183 a_n1451_2298# a_n1551_2201# a_n1609_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X184 a_1551_2298# a_1451_2201# a_1393_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X185 a_n503_1426# a_n603_1329# a_n661_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X186 a_n1293_n1190# a_n1393_n1287# a_n1451_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X187 a_129_1862# a_29_1765# a_n29_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X188 a_n345_554# a_n445_457# a_n503_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X189 a_n1135_n2498# a_n1235_n2595# a_n1293_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X190 a_n187_n1626# a_n287_n1723# a_n345_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X191 a_1551_n2934# a_1451_n3031# a_1393_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X192 a_n29_n2934# a_n129_n3031# a_n187_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X193 a_n503_n2062# a_n603_n2159# a_n661_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X194 a_n977_2734# a_n1077_2637# a_n1135_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X195 a_1551_n1190# a_1451_n1287# a_1393_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X196 a_n29_n1190# a_n129_n1287# a_n187_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X197 a_1077_118# a_977_21# a_919_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X198 a_445_1862# a_345_1765# a_287_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X199 a_287_n2062# a_187_n2159# a_129_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X200 a_1077_2734# a_977_2637# a_919_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X201 a_n503_2734# a_n603_2637# a_n661_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X202 a_n345_n754# a_n445_n851# a_n503_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X203 a_n1293_n2498# a_n1393_n2595# a_n1451_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X204 a_1551_1862# a_1451_1765# a_1393_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X205 a_n661_990# a_n761_893# a_n819_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X206 a_1551_118# a_1451_21# a_1393_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X207 a_n977_n318# a_n1077_n415# a_n1135_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X208 a_n187_n2934# a_n287_n3031# a_n345_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X209 a_n1451_1862# a_n1551_1765# a_n1609_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X210 a_n29_n2498# a_n129_n2595# a_n187_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X211 a_n661_n2062# a_n761_n2159# a_n819_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X212 a_n187_n1190# a_n287_n1287# a_n345_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X213 a_n977_2298# a_n1077_2201# a_n1135_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X214 a_n503_554# a_n603_457# a_n661_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X215 a_1551_n2498# a_1451_n2595# a_1393_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X216 a_n29_1426# a_n129_1329# a_n187_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X217 a_603_1426# a_503_1329# a_445_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X218 a_129_990# a_29_893# a_n29_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X219 a_1077_n318# a_977_n415# a_919_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X220 a_1077_2298# a_977_2201# a_919_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X221 a_n503_n318# a_n603_n415# a_n661_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X222 a_129_n754# a_29_n851# a_n29_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X223 a_n503_2298# a_n603_2201# a_n661_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X224 a_n187_990# a_n287_893# a_n345_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X225 a_761_118# a_661_21# a_603_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X226 a_n187_n2498# a_n287_n2595# a_n345_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X227 a_n1135_n2062# a_n1235_n2159# a_n1293_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X228 a_129_n1626# a_29_n1723# a_n29_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X229 a_n29_2734# a_n129_2637# a_n187_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X230 a_603_2734# a_503_2637# a_445_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X231 a_n29_554# a_n129_457# a_n187_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X232 a_445_n754# a_345_n851# a_287_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X233 a_n977_1862# a_n1077_1765# a_n1135_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X234 a_n1451_n754# a_n1551_n851# a_n1609_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X235 a_1551_n754# a_1451_n851# a_1393_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X236 a_1077_1862# a_977_1765# a_919_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X237 a_n819_990# a_n919_893# a_n977_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X238 a_287_118# a_187_21# a_129_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X239 a_n1293_n2062# a_n1393_n2159# a_n1451_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X240 a_n503_1862# a_n603_1765# a_n661_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X241 a_1393_554# a_1293_457# a_1235_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X242 a_n29_n318# a_n129_n415# a_n187_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X243 a_603_n318# a_503_n415# a_445_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X244 a_129_n2934# a_29_n3031# a_n29_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X245 a_1235_1426# a_1135_1329# a_1077_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X246 a_n345_990# a_n445_893# a_n503_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X247 a_1235_118# a_1135_21# a_1077_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X248 a_129_n1190# a_29_n1287# a_n29_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X249 a_n29_2298# a_n129_2201# a_n187_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X250 a_603_2298# a_503_2201# a_445_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X251 a_n1135_1426# a_n1235_1329# a_n1293_1426# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X252 a_1551_n2062# a_1451_n2159# a_1393_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X253 a_n29_n2062# a_n129_n2159# a_n187_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X254 a_445_n1626# a_345_n1723# a_287_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X255 a_1077_554# a_977_457# a_919_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X256 a_919_118# a_819_21# a_761_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X257 a_n1135_2734# a_n1235_2637# a_n1293_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X258 a_1235_2734# a_1135_2637# a_1077_2734# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X259 a_1551_554# a_1451_457# a_1393_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X260 a_445_118# a_345_21# a_287_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X261 a_129_n2498# a_29_n2595# a_n29_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X262 a_n187_n2062# a_n287_n2159# a_n345_n2062# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X263 a_n977_n754# a_n1077_n851# a_n1135_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X264 a_445_n2934# a_345_n3031# a_287_n2934# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X265 a_n503_990# a_n603_893# a_n661_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X266 a_445_n1190# a_345_n1287# a_287_n1190# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X267 a_n29_1862# a_n129_1765# a_n187_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X268 a_603_1862# a_503_1765# a_445_1862# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X269 a_1077_n754# a_977_n851# a_919_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X270 a_1235_n318# a_1135_n415# a_1077_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X271 a_n503_n754# a_n603_n851# a_n661_n754# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X272 a_919_n1626# a_819_n1723# a_761_n1626# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X273 a_n1135_n318# a_n1235_n415# a_n1293_n318# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X274 a_1235_2298# a_1135_2201# a_1077_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X275 a_761_554# a_661_457# a_603_554# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X276 a_n1135_2298# a_n1235_2201# a_n1293_2298# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X277 a_603_118# a_503_21# a_445_118# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X278 a_n29_990# a_n129_893# a_n187_990# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X279 a_445_n2498# a_345_n2595# a_287_n2498# w_n1809_n3231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_H7BQFY a_n287_n188# a_n29_n100# a_n187_n100#
+ a_n345_n100# a_129_n100# a_287_n100# a_n479_n322# a_29_n188# a_n129_n188# a_187_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n187_n100# a_n287_n188# a_n345_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X2 a_n29_n100# a_n129_n188# a_n187_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_287_n100# a_187_n188# a_129_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_H7BQ24 a_n287_n188# a_n29_n100# a_n187_n100#
+ a_n345_n100# a_129_n100# a_287_n100# a_n479_n322# a_29_n188# a_n129_n188# a_187_n188#
X0 a_129_n100# a_29_n188# a_n29_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 a_n187_n100# a_n287_n188# a_n345_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X2 a_n29_n100# a_n129_n188# a_n187_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 a_287_n100# a_187_n188# a_129_n100# a_n479_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

.subckt follower_amp vdd out ena in vsub vss
XXM12 m1_651_3930# m1_651_3930# out m1_651_3930# vdd out vdd m1_651_3930# vdd out
+ vdd out out m1_651_3930# out vdd m1_651_3930# m1_651_3930# vdd vdd out m1_651_3930#
+ m1_651_3930# out m1_651_3930# m1_651_3930# out vdd m1_651_3930# m1_651_3930# m1_651_3930#
+ out m1_651_3930# m1_651_3930# vdd vdd vdd m1_651_3930# m1_651_3930# m1_651_3930#
+ m1_651_3930# out sky130_fd_pr__pfet_g5v0d10v5_AQ2WAW
XXM13 m1_2399_1244# vss nbias ena sky130_fd_pr__nfet_g5v0d10v5_UNEQFS
XXM24 pbias vss vss nbias sky130_fd_pr__nfet_g5v0d10v5_UNEQFS
XXM25 pbias vdd pbias vcomp vdd vdd pbias pbias sky130_fd_pr__pfet_g5v0d10v5_KLJMY6
XXM27 vcomp m2_526_2596# vdd vcomp out in out m1_811_2614# in vcomp sky130_fd_pr__pfet_g5v0d10v5_KLWMS5
XXM29 m1_811_2614# vss vss m1_811_2614# sky130_fd_pr__nfet_g5v0d10v5_UNEQFS
XXR1 m1_3337_606# vdd m1_604_772# m1_604_772# m1_2399_1244# m1_3337_606# vss sky130_fd_pr__res_xhigh_po_0p35_HLA228
XXM1 vss m2_1742_2323# m1_505_3709# m2_1930_2454# out in sky130_fd_pr__nfet_g5v0d10v5_FJGQFC
XXM5 vdd m1_505_3709# vdd vdd m2_1930_2454# m2_1930_2454# m2_1930_2454# m2_1930_2454#
+ m2_1930_2454# vdd sky130_fd_pr__pfet_g5v0d10v5_KLWMS5
XXXD1 vss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__0
XXM6 vdd m1_651_3930# vdd vdd m2_3105_2460# m2_3105_2460# m2_3105_2460# m2_3105_2460#
+ m2_3105_2460# vdd sky130_fd_pr__pfet_g5v0d10v5_KLWMS5
XXXD2 vss in sky130_fd_pr__diode_pw2nd_05v5_FT76RJ__0
XXM7 vss vss m2_2845_2323# m2_2845_2323# nbias nbias sky130_fd_pr__nfet_g5v0d10v5_XJGQ2Y
XXM8 vss vss m2_1742_2323# nbias sky130_fd_pr__nfet_g5v0d10v5_UNEQFS
XXM9 m2_2845_2323# m2_3105_2460# in vss m1_651_3930# out sky130_fd_pr__nfet_05v0_nvt_BH6ZTK
XXM30 m2_526_2596# vss vss m1_811_2614# sky130_fd_pr__nfet_g5v0d10v5_UNEQFS
XXM20 out vdd m1_505_3709# out vdd out m1_505_3709# out m1_505_3709# m1_505_3709#
+ vdd m1_505_3709# m1_505_3709# vdd m1_505_3709# out vdd m1_505_3709# out m1_505_3709#
+ out out m1_505_3709# m1_505_3709# m1_505_3709# vdd vdd out out m1_505_3709# vdd
+ m1_505_3709# m1_505_3709# vdd out vdd m1_505_3709# m1_505_3709# m1_505_3709# vdd
+ out out m1_505_3709# vdd vdd m1_505_3709# m1_505_3709# m1_505_3709# out m1_505_3709#
+ vdd m1_505_3709# m1_505_3709# vdd out m1_505_3709# m1_505_3709# m1_505_3709# vdd
+ vdd out vdd m1_505_3709# m1_505_3709# vdd out vdd m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# out out out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# out
+ m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709#
+ vdd m1_505_3709# out out out m1_505_3709# m1_505_3709# out vdd m1_505_3709# m1_505_3709#
+ out m1_505_3709# out m1_505_3709# vdd out m1_505_3709# vdd out vdd m1_505_3709#
+ out m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709# vdd vdd m1_505_3709#
+ vdd m1_505_3709# vdd m1_505_3709# out m1_505_3709# out out m1_505_3709# vdd out
+ out out m1_505_3709# vdd vdd m1_505_3709# vdd m1_505_3709# out m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# out m1_505_3709# vdd vdd m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# vdd m1_505_3709# m1_505_3709# out m1_505_3709# vdd m1_505_3709# out
+ m1_505_3709# m1_505_3709# out m1_505_3709# vdd out m1_505_3709# vdd m1_505_3709#
+ vdd m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709# out vdd m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# vdd out vdd
+ vdd m1_505_3709# out out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709#
+ out m1_505_3709# out m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ out vdd m1_505_3709# m1_505_3709# m1_505_3709# vdd out out m1_505_3709# m1_505_3709#
+ out vdd m1_505_3709# m1_505_3709# out m1_505_3709# out vdd m1_505_3709# m1_505_3709#
+ m1_505_3709# out out vdd out m1_505_3709# out vdd m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# vdd m1_505_3709# out out vdd vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ vdd out m1_505_3709# m1_505_3709# out m1_505_3709# out m1_505_3709# m1_505_3709#
+ vdd out m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# m1_505_3709# vdd
+ out m1_505_3709# out m1_505_3709# m1_505_3709# vdd out out vdd m1_505_3709# m1_505_3709#
+ out out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# out out m1_505_3709#
+ vdd m1_505_3709# m1_505_3709# m1_505_3709# out m1_505_3709# m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# m1_505_3709# out vdd m1_505_3709# vdd m1_505_3709# vdd out vdd out
+ out m1_505_3709# vdd vdd out out out m1_505_3709# m1_505_3709# m1_505_3709# out
+ out vdd out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# vdd out out vdd m1_505_3709# m1_505_3709# m1_505_3709#
+ out m1_505_3709# m1_505_3709# m1_505_3709# vdd vdd vdd out vdd m1_505_3709# vdd
+ out out m1_505_3709# out m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709#
+ m1_505_3709# vdd m1_505_3709# m1_505_3709# vdd vdd m1_505_3709# m1_505_3709# vdd
+ out m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# vdd vdd out vdd m1_505_3709#
+ m1_505_3709# vdd out vdd out m1_505_3709# out m1_505_3709# out m1_505_3709# out
+ m1_505_3709# vdd m1_505_3709# out m1_505_3709# vdd out out vdd m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# out vdd vdd m1_505_3709# m1_505_3709# out vdd vdd vdd
+ vdd m1_505_3709# vdd m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709#
+ out vdd m1_505_3709# out vdd out out m1_505_3709# out out m1_505_3709# vdd m1_505_3709#
+ vdd m1_505_3709# vdd out vdd m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# vdd m1_505_3709# m1_505_3709# vdd m1_505_3709#
+ vdd out m1_505_3709# m1_505_3709# vdd out vdd out m1_505_3709# vdd out m1_505_3709#
+ m1_505_3709# vdd m1_505_3709# vdd m1_505_3709# out m1_505_3709# out vdd out vdd
+ out m1_505_3709# m1_505_3709# vdd vdd out out m1_505_3709# out m1_505_3709# m1_505_3709#
+ out m1_505_3709# m1_505_3709# vdd out out m1_505_3709# vdd vdd out out vdd m1_505_3709#
+ out m1_505_3709# vdd out m1_505_3709# m1_505_3709# vdd out m1_505_3709# vdd m1_505_3709#
+ m1_505_3709# m1_505_3709# m1_505_3709# m1_505_3709# out out out vdd m1_505_3709#
+ vdd out m1_505_3709# out vdd out m1_505_3709# vdd out out vdd out m1_505_3709# m1_505_3709#
+ vdd out m1_505_3709# out vdd vdd out vdd out out m1_505_3709# vdd m1_505_3709# vdd
+ m1_505_3709# m1_505_3709# m1_505_3709# out out m1_505_3709# m1_505_3709# vdd out
+ m1_505_3709# m1_505_3709# out sky130_fd_pr__pfet_g5v0d10v5_Z8JNCQ
XXM10 nbias vss nbias vss nbias vss vss nbias nbias nbias sky130_fd_pr__nfet_g5v0d10v5_H7BQFY
XXM22 m2_526_2596# vss out vss out vss vss m2_526_2596# m2_526_2596# m2_526_2596#
+ sky130_fd_pr__nfet_g5v0d10v5_H7BQ24
.ends

.subckt dac_3v_column b4b dum1_out b0_uq12 b0_uq1 b2b_uq0 dac_3v_cell_top_0/m4_97_801#
+ b0_uq11 b0_uq10 b2b_uq2 b3b b4 b0b_uq13 b2b_uq1 b0_uq6 dac_3v_cell_0[2]/w_316_892#
+ dum0_in dac_3v_cell_0[1]/w_316_892# b0b_uq11 b0 dac_3v_cell_top_0/m4_97_1059# b1
+ b0b_uq10 b1_uq6 dac_3v_cell_0[6]/w_316_892# b0b_uq12 b1_uq1 b1_uq2 b1_uq0 b3 b0_uq3
+ b0b_uq2 b1_uq3 b0b_uq1 b0_uq14 dac_3v_cell_0[5]/w_316_892# b0b_uq14 b0b_uq7 b0b_uq0
+ b0_uq2 b0b_uq6 out_5 b0b_uq9 out_4 dac_3v_cell_top_0/m1_290_591# b0b_uq8 b1b_uq6
+ b0_uq13 b3_uq0 b3b_uq0 b1b_uq5 dac_3v_cell_0[4]/w_316_892# b2_uq1 res0_in b2 m2_801_196#
+ b1b_uq4 b0_uq5 b0_uq0 b2_uq0 b1b_uq3 b0_uq4 b1b_uq2 b1_uq5 b2_uq2 m2_791_1314# b1_uq4
+ b1b_uq0 b0b_uq5 m2_791_14877# dac_3v_cell_0[7]/w_316_892# b0_uq9 b0b b1b_uq1 res1_out
+ dac_3v_cell_top_0/m1_290_1114# b0_uq8 dac_3v_cell_0[3]/w_316_892# b1b b0b_uq4 b0b_uq3
+ b0_uq7 m2_801_13759# b2b VSUBS
Xdac_3v_cell_0[0] m2_791_1314# m2_801_196# m2_328_1119# m2_328_1119# res1_out m2_791_1314#
+ VSUBS m2_449_485# m2_328_1119# dum1_out m2_801_196# m2_449_485# VSUBS m2_449_485#
+ VSUBS m2_791_1314# m2_801_196# VSUBS res0_in dum0_in VSUBS dac_3v_cell
Xdac_3v_cell_0[1] b0b m2_791_1314# out0_0_0 out0_1_0 dac_3v_cell_0[1]/m1_824_799#
+ b1b_uq0 VSUBS out0_0_0 out1_0_3 res1_out b0_uq0 out_3 b4b out_4 b0 dac_3v_cell_0[1]/w_316_892#
+ b4 b1_uq0 dac_3v_cell_0[2]/m1_155_n223# res0_in b0b_uq0 dac_3v_cell
Xdac_3v_cell_0[2] b0_uq2 dac_3v_cell_0[1]/w_316_892# out0_2 out0_1_0 dac_3v_cell_0[2]/m1_824_799#
+ b2b_uq0 VSUBS out0_0_0 out1_0_3 dac_3v_cell_0[1]/m1_824_799# b0b_uq1 out1_1_1 b1b
+ out1_0_3 b0b_uq2 dac_3v_cell_0[2]/w_316_892# b1 b2_uq0 dac_3v_cell_0[3]/m1_155_n223#
+ dac_3v_cell_0[2]/m1_155_n223# b0_uq1 dac_3v_cell
Xdac_3v_cell_0[3] b0b_uq4 dac_3v_cell_0[2]/w_316_892# out0_0_1 out0_1_0 dac_3v_cell_0[3]/m1_824_799#
+ b1_uq1 VSUBS out0_0_1 out1_0_2 dac_3v_cell_0[2]/m1_824_799# b0_uq3 out1_1_1 b2b
+ out1_2 b0_uq4 dac_3v_cell_0[3]/w_316_892# b2 b1b_uq1 dac_3v_cell_0[4]/m1_155_n223#
+ dac_3v_cell_0[3]/m1_155_n223# b0b_uq3 dac_3v_cell
Xdac_3v_cell_0[4] b0_uq6 dac_3v_cell_0[3]/w_316_892# out_3 out0_2 dac_3v_cell_0[4]/m1_824_799#
+ b3b_uq0 VSUBS out0_0_1 out1_0_2 dac_3v_cell_0[3]/m1_824_799# b0b_uq5 out1_1_1 b1_uq2
+ out1_0_2 b0b_uq6 dac_3v_cell_0[4]/w_316_892# b1b_uq2 b3_uq0 dac_3v_cell_0[5]/m1_155_n223#
+ dac_3v_cell_0[4]/m1_155_n223# b0_uq5 dac_3v_cell
Xdac_3v_cell_0[5] b0b_uq8 dac_3v_cell_0[4]/w_316_892# out0_0_2 out0_1_1 dac_3v_cell_0[5]/m1_824_799#
+ b1b_uq3 VSUBS out0_0_2 out1_0_1 dac_3v_cell_0[4]/m1_824_799# b0_uq7 out1_2 b3b out_3
+ b0_uq8 dac_3v_cell_0[5]/w_316_892# b3 b1_uq3 dac_3v_cell_0[6]/m1_155_n223# dac_3v_cell_0[5]/m1_155_n223#
+ b0b_uq7 dac_3v_cell
Xdac_3v_cell_0[6] b0_uq10 dac_3v_cell_0[5]/w_316_892# out0_2 out0_1_1 dac_3v_cell_0[6]/m1_824_799#
+ b2_uq1 VSUBS out0_0_2 out1_0_1 dac_3v_cell_0[5]/m1_824_799# b0b_uq9 out1_1_0 b1b_uq4
+ out1_0_1 b0b_uq10 dac_3v_cell_0[6]/w_316_892# b1_uq4 b2b_uq1 dac_3v_cell_0[7]/m1_155_n223#
+ dac_3v_cell_0[6]/m1_155_n223# b0_uq9 dac_3v_cell
Xdac_3v_cell_0[7] b0b_uq12 dac_3v_cell_0[6]/w_316_892# out0_0_3 out0_1_1 dac_3v_cell_0[7]/m1_824_799#
+ b1_uq5 VSUBS out0_0_3 out1_0_0 dac_3v_cell_0[6]/m1_824_799# b0_uq11 out1_1_0 b2_uq2
+ out1_2 b0_uq12 dac_3v_cell_0[7]/w_316_892# b2b_uq2 b1b_uq5 dac_3v_cell_top_0/m1_155_n223#
+ dac_3v_cell_0[7]/m1_155_n223# b0b_uq11 dac_3v_cell
Xdac_3v_cell_1 m2_791_14877# m2_801_13759# m2_330_14682# m2_330_14682# dum0_out m2_791_14877#
+ VSUBS m2_449_14048# m2_330_14682# res1_in m2_801_13759# m2_449_14048# VSUBS m2_449_14048#
+ VSUBS m2_791_14877# m2_801_13759# VSUBS dum0_out res1_in VSUBS dac_3v_cell
Xdac_3v_cell_top_0 b0_uq14 dac_3v_cell_0[7]/w_316_892# out_4 out_5 res1_in m2_801_13759#
+ dac_3v_cell_top_0/m1_290_1114# VSUBS out0_0_3 out1_0_0 dac_3v_cell_0[7]/m1_824_799#
+ b0b_uq13 dac_3v_cell_top_0/m4_97_801# out1_1_0 dac_3v_cell_top_0/m4_97_1059# b1_uq6
+ out1_0_0 b0b_uq14 b1b_uq6 dac_3v_cell_top_0/m1_290_591# dac_3v_cell_top_0/m1_155_n223#
+ b0_uq13 dac_3v_cell_top
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_4AXGXB__0 a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt rdac_level_shifter dvdd bitb_out bit_out bit_in avdd agnd
Xsky130_fd_sc_hvl__inv_8_1 bitb_out agnd agnd avdd avdd bit_out sky130_fd_sc_hvl__inv_8
Xsky130_fd_sc_hvl__inv_4_0 sky130_fd_sc_hvl__inv_4_0/A agnd agnd avdd avdd sky130_fd_sc_hvl__inv_8_0/A
+ sky130_fd_sc_hvl__inv_4
Xsky130_fd_sc_hvl__inv_2_0 sky130_fd_sc_hvl__inv_2_0/A agnd agnd avdd avdd sky130_fd_sc_hvl__inv_4_0/A
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0 bit_in dvdd agnd avdd avdd sky130_fd_sc_hvl__inv_2_0/A
+ avdd agnd agnd sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_pr__diode_pw2nd_05v5_4AXGXB_0 agnd bit_in sky130_fd_pr__diode_pw2nd_05v5_4AXGXB__0
Xsky130_fd_sc_hvl__inv_8_0 sky130_fd_sc_hvl__inv_8_0/A agnd agnd avdd avdd bitb_out
+ sky130_fd_sc_hvl__inv_8
.ends

.subckt level_shifter_array rdac_level_shifter_0[2]/bit_out rdac_level_shifter_0[6]/bitb_out
+ rdac_level_shifter_0[2]/bitb_out rdac_level_shifter_0[3]/bit_in rdac_level_shifter_0[7]/bit_in
+ rdac_level_shifter_0[6]/bit_out rdac_level_shifter_0[3]/bit_out rdac_level_shifter_0[7]/dvdd
+ rdac_level_shifter_0[0]/bit_in rdac_level_shifter_0[3]/bitb_out rdac_level_shifter_0[0]/bit_out
+ rdac_level_shifter_0[4]/bit_in rdac_level_shifter_0[7]/bit_out rdac_level_shifter_0[4]/bit_out
+ rdac_level_shifter_0[4]/bitb_out rdac_level_shifter_0[1]/bit_in rdac_level_shifter_0[0]/bitb_out
+ rdac_level_shifter_0[5]/bit_in rdac_level_shifter_0[1]/bit_out rdac_level_shifter_0[7]/bitb_out
+ rdac_level_shifter_0[5]/bitb_out rdac_level_shifter_0[5]/bit_out rdac_level_shifter_0[2]/bit_in
+ rdac_level_shifter_0[1]/bitb_out VSUBS rdac_level_shifter_0[6]/bit_in rdac_level_shifter_0[7]/avdd
Xrdac_level_shifter_0[0] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[0]/bitb_out
+ rdac_level_shifter_0[0]/bit_out rdac_level_shifter_0[0]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
Xrdac_level_shifter_0[1] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[1]/bitb_out
+ rdac_level_shifter_0[1]/bit_out rdac_level_shifter_0[1]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
Xrdac_level_shifter_0[2] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[2]/bitb_out
+ rdac_level_shifter_0[2]/bit_out rdac_level_shifter_0[2]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
Xrdac_level_shifter_0[3] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[3]/bitb_out
+ rdac_level_shifter_0[3]/bit_out rdac_level_shifter_0[3]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
Xrdac_level_shifter_0[4] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[4]/bitb_out
+ rdac_level_shifter_0[4]/bit_out rdac_level_shifter_0[4]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
Xrdac_level_shifter_0[5] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[5]/bitb_out
+ rdac_level_shifter_0[5]/bit_out rdac_level_shifter_0[5]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
Xrdac_level_shifter_0[6] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[6]/bitb_out
+ rdac_level_shifter_0[6]/bit_out rdac_level_shifter_0[6]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
Xrdac_level_shifter_0[7] rdac_level_shifter_0[7]/dvdd rdac_level_shifter_0[7]/bitb_out
+ rdac_level_shifter_0[7]/bit_out rdac_level_shifter_0[7]/bit_in rdac_level_shifter_0[7]/avdd
+ VSUBS rdac_level_shifter
.ends

.subckt dac_3v_cell_dummy m4_99_18# w_318_n275# m4_99_276# m4_99_801# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ m4_99_930# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732# m4_99_405# m4_99_1059#
+ m4_99_672# w_316_892# sky130_fd_pr__res_high_po_0p35_AW5QUD_0/a_n35_300# m4_99_147#
+ m1_155_n223# m1_824_799#
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_0 sky130_fd_pr__res_high_po_0p35_AW5QUD_0/a_n35_300#
+ m1_155_n223# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__res_high_po_0p35_AW5QUD_1 m1_824_799# sky130_fd_pr__res_high_po_0p35_AW5QUD_1/a_n35_n732#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__res_high_po_0p35_AW5QUD
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_0 m1_387_847# m1_387_847# w_316_892# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_1 m1_824_799# m1_387_847# w_316_892# w_316_892#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_2 m1_545_212# m1_545_212# w_318_n275# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__pfet_g5v0d10v5_9992MR_3 m1_545_212# m1_155_n223# w_318_n275# w_318_n275#
+ sky130_fd_pr__pfet_g5v0d10v5_9992MR__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_0 m1_387_847# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ m1_387_847# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_1 m1_387_847# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ m1_824_799# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_2 m1_155_n223# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ m1_545_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
Xsky130_fd_pr__nfet_g5v0d10v5_NHLDUY_3 m1_545_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS
+ m1_545_212# sky130_fd_pr__pfet_g5v0d10v5_9992MR_3/VSUBS sky130_fd_pr__nfet_g5v0d10v5_NHLDUY__0
.ends

.subckt dac_3v_column_dummy m1_988_1608# dac_3v_cell_dummy_0[6]/m4_99_147# dac_3v_cell_dummy_0[0]/w_318_n275#
+ dac_3v_cell_dummy_0[7]/m4_99_147# dac_3v_cell_dummy_0[6]/m4_99_18# dac_3v_cell_dummy_0[8]/m4_99_147#
+ dac_3v_cell_dummy_0[9]/m4_99_147# dac_3v_cell_dummy_0[7]/m4_99_18# dac_3v_cell_dummy_0[0]/m4_99_276#
+ dac_3v_cell_dummy_0[0]/m4_99_801# dac_3v_cell_dummy_0[1]/m4_99_276# dac_3v_cell_dummy_0[7]/m4_99_1059#
+ dac_3v_cell_dummy_0[2]/m4_99_1059# dac_3v_cell_dummy_0[1]/m4_99_801# dac_3v_cell_dummy_0[2]/m4_99_276#
+ dac_3v_cell_dummy_0[2]/m4_99_801# dac_3v_cell_dummy_0[3]/m4_99_276# dac_3v_cell_dummy_0[3]/m4_99_801#
+ dac_3v_cell_dummy_0[4]/m4_99_276# dac_3v_cell_dummy_0[8]/m4_99_18# dac_3v_cell_dummy_0[4]/m4_99_801#
+ dac_3v_cell_dummy_0[5]/m4_99_276# dac_3v_cell_dummy_0[5]/m4_99_801# dac_3v_cell_dummy_0[6]/m4_99_276#
+ dac_3v_cell_dummy_0[6]/m4_99_801# dac_3v_cell_dummy_0[7]/m4_99_276# dac_3v_cell_dummy_0[7]/m4_99_801#
+ dac_3v_cell_dummy_0[9]/m4_99_18# dac_3v_cell_dummy_0[8]/m4_99_276# dac_3v_cell_dummy_0[8]/m4_99_801#
+ dac_3v_cell_dummy_0[9]/m4_99_276# dac_3v_cell_dummy_0[9]/m4_99_801# dac_3v_cell_dummy_0[6]/m4_99_1059#
+ dac_3v_cell_dummy_0[1]/m4_99_1059# dac_3v_cell_dummy_0[0]/m4_99_930# dac_3v_cell_dummy_0[1]/m4_99_930#
+ dac_3v_cell_dummy_0[2]/m4_99_930# dac_3v_cell_dummy_0[3]/m4_99_930# dac_3v_cell_dummy_0[0]/m4_99_18#
+ dac_3v_cell_dummy_0[4]/m4_99_930# dac_3v_cell_dummy_0[5]/m4_99_930# dac_3v_cell_dummy_0[6]/m4_99_930#
+ VSUBS dac_3v_cell_dummy_0[5]/m4_99_1059# dac_3v_cell_dummy_0[7]/m4_99_930# dac_3v_cell_dummy_0[1]/m4_99_18#
+ dac_3v_cell_dummy_0[0]/m4_99_1059# dac_3v_cell_dummy_0[8]/m4_99_930# dac_3v_cell_dummy_0[9]/m4_99_930#
+ dac_3v_cell_dummy_0[0]/m4_99_405# dac_3v_cell_dummy_0[1]/m4_99_405# dac_3v_cell_dummy_0[2]/m4_99_405#
+ dac_3v_cell_dummy_0[0]/m4_99_672# dac_3v_cell_dummy_0[2]/m4_99_18# dac_3v_cell_dummy_0[3]/m4_99_405#
+ m1_938_45# dac_3v_cell_dummy_0[1]/m4_99_672# dac_3v_cell_dummy_0[4]/m4_99_405# dac_3v_cell_dummy_0[2]/m4_99_672#
+ dac_3v_cell_dummy_0[1]/w_316_892# dac_3v_cell_dummy_0[5]/m4_99_405# dac_3v_cell_dummy_0[3]/m4_99_672#
+ dac_3v_cell_dummy_0[2]/w_316_892# dac_3v_cell_dummy_0[4]/m4_99_672# dac_3v_cell_dummy_0[6]/m4_99_405#
+ dac_3v_cell_dummy_0[9]/m4_99_1059# dac_3v_cell_dummy_0[3]/m4_99_18# dac_3v_cell_dummy_0[4]/m4_99_1059#
+ dac_3v_cell_dummy_0[3]/w_316_892# dac_3v_cell_dummy_0[5]/m4_99_672# dac_3v_cell_dummy_0[7]/m4_99_405#
+ dac_3v_cell_dummy_0[8]/m4_99_405# dac_3v_cell_dummy_0[6]/m4_99_672# dac_3v_cell_dummy_0[4]/w_316_892#
+ dac_3v_cell_dummy_0[0]/w_316_892# dac_3v_cell_dummy_0[7]/m4_99_672# dac_3v_cell_dummy_0[9]/m4_99_405#
+ dac_3v_cell_dummy_0[5]/w_316_892# dac_3v_cell_dummy_0[6]/w_316_892# dac_3v_cell_dummy_0[8]/m4_99_672#
+ dac_3v_cell_dummy_0[4]/m4_99_18# dac_3v_cell_dummy_0[7]/w_316_892# dac_3v_cell_dummy_0[0]/m4_99_147#
+ dac_3v_cell_dummy_0[9]/m4_99_672# dac_3v_cell_dummy_0[8]/w_316_892# dac_3v_cell_dummy_0[1]/m4_99_147#
+ m1_n18_1607# dac_3v_cell_dummy_0[9]/w_316_892# dac_3v_cell_dummy_0[2]/m4_99_147#
+ dac_3v_cell_dummy_0[3]/m4_99_147# dac_3v_cell_dummy_0[5]/m4_99_18# m1_n18_45# dac_3v_cell_dummy_0[8]/m4_99_1059#
+ dac_3v_cell_dummy_0[4]/m4_99_147# dac_3v_cell_dummy_0[3]/m4_99_1059# dac_3v_cell_dummy_0[5]/m4_99_147#
Xdac_3v_cell_dummy_0[0] dac_3v_cell_dummy_0[0]/m4_99_18# dac_3v_cell_dummy_0[0]/w_318_n275#
+ dac_3v_cell_dummy_0[0]/m4_99_276# dac_3v_cell_dummy_0[0]/m4_99_801# VSUBS dac_3v_cell_dummy_0[0]/m4_99_930#
+ m1_938_45# dac_3v_cell_dummy_0[0]/m4_99_405# dac_3v_cell_dummy_0[0]/m4_99_1059#
+ dac_3v_cell_dummy_0[0]/m4_99_672# dac_3v_cell_dummy_0[0]/w_316_892# m1_n18_1607#
+ dac_3v_cell_dummy_0[0]/m4_99_147# m1_n18_45# m1_988_1608# dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[1] dac_3v_cell_dummy_0[1]/m4_99_18# dac_3v_cell_dummy_0[0]/w_316_892#
+ dac_3v_cell_dummy_0[1]/m4_99_276# dac_3v_cell_dummy_0[1]/m4_99_801# VSUBS dac_3v_cell_dummy_0[1]/m4_99_930#
+ m1_988_1608# dac_3v_cell_dummy_0[1]/m4_99_405# dac_3v_cell_dummy_0[1]/m4_99_1059#
+ dac_3v_cell_dummy_0[1]/m4_99_672# dac_3v_cell_dummy_0[1]/w_316_892# dac_3v_cell_dummy_0[2]/m1_155_n223#
+ dac_3v_cell_dummy_0[1]/m4_99_147# m1_n18_1607# dac_3v_cell_dummy_0[1]/m1_824_799#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[2] dac_3v_cell_dummy_0[2]/m4_99_18# dac_3v_cell_dummy_0[1]/w_316_892#
+ dac_3v_cell_dummy_0[2]/m4_99_276# dac_3v_cell_dummy_0[2]/m4_99_801# VSUBS dac_3v_cell_dummy_0[2]/m4_99_930#
+ dac_3v_cell_dummy_0[1]/m1_824_799# dac_3v_cell_dummy_0[2]/m4_99_405# dac_3v_cell_dummy_0[2]/m4_99_1059#
+ dac_3v_cell_dummy_0[2]/m4_99_672# dac_3v_cell_dummy_0[2]/w_316_892# dac_3v_cell_dummy_0[3]/m1_155_n223#
+ dac_3v_cell_dummy_0[2]/m4_99_147# dac_3v_cell_dummy_0[2]/m1_155_n223# dac_3v_cell_dummy_0[2]/m1_824_799#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[3] dac_3v_cell_dummy_0[3]/m4_99_18# dac_3v_cell_dummy_0[2]/w_316_892#
+ dac_3v_cell_dummy_0[3]/m4_99_276# dac_3v_cell_dummy_0[3]/m4_99_801# VSUBS dac_3v_cell_dummy_0[3]/m4_99_930#
+ dac_3v_cell_dummy_0[2]/m1_824_799# dac_3v_cell_dummy_0[3]/m4_99_405# dac_3v_cell_dummy_0[3]/m4_99_1059#
+ dac_3v_cell_dummy_0[3]/m4_99_672# dac_3v_cell_dummy_0[3]/w_316_892# dac_3v_cell_dummy_0[4]/m1_155_n223#
+ dac_3v_cell_dummy_0[3]/m4_99_147# dac_3v_cell_dummy_0[3]/m1_155_n223# dac_3v_cell_dummy_0[3]/m1_824_799#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[4] dac_3v_cell_dummy_0[4]/m4_99_18# dac_3v_cell_dummy_0[3]/w_316_892#
+ dac_3v_cell_dummy_0[4]/m4_99_276# dac_3v_cell_dummy_0[4]/m4_99_801# VSUBS dac_3v_cell_dummy_0[4]/m4_99_930#
+ dac_3v_cell_dummy_0[3]/m1_824_799# dac_3v_cell_dummy_0[4]/m4_99_405# dac_3v_cell_dummy_0[4]/m4_99_1059#
+ dac_3v_cell_dummy_0[4]/m4_99_672# dac_3v_cell_dummy_0[4]/w_316_892# dac_3v_cell_dummy_0[5]/m1_155_n223#
+ dac_3v_cell_dummy_0[4]/m4_99_147# dac_3v_cell_dummy_0[4]/m1_155_n223# dac_3v_cell_dummy_0[4]/m1_824_799#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[5] dac_3v_cell_dummy_0[5]/m4_99_18# dac_3v_cell_dummy_0[4]/w_316_892#
+ dac_3v_cell_dummy_0[5]/m4_99_276# dac_3v_cell_dummy_0[5]/m4_99_801# VSUBS dac_3v_cell_dummy_0[5]/m4_99_930#
+ dac_3v_cell_dummy_0[4]/m1_824_799# dac_3v_cell_dummy_0[5]/m4_99_405# dac_3v_cell_dummy_0[5]/m4_99_1059#
+ dac_3v_cell_dummy_0[5]/m4_99_672# dac_3v_cell_dummy_0[5]/w_316_892# dac_3v_cell_dummy_0[6]/m1_155_n223#
+ dac_3v_cell_dummy_0[5]/m4_99_147# dac_3v_cell_dummy_0[5]/m1_155_n223# dac_3v_cell_dummy_0[5]/m1_824_799#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[6] dac_3v_cell_dummy_0[6]/m4_99_18# dac_3v_cell_dummy_0[5]/w_316_892#
+ dac_3v_cell_dummy_0[6]/m4_99_276# dac_3v_cell_dummy_0[6]/m4_99_801# VSUBS dac_3v_cell_dummy_0[6]/m4_99_930#
+ dac_3v_cell_dummy_0[5]/m1_824_799# dac_3v_cell_dummy_0[6]/m4_99_405# dac_3v_cell_dummy_0[6]/m4_99_1059#
+ dac_3v_cell_dummy_0[6]/m4_99_672# dac_3v_cell_dummy_0[6]/w_316_892# dac_3v_cell_dummy_0[7]/m1_155_n223#
+ dac_3v_cell_dummy_0[6]/m4_99_147# dac_3v_cell_dummy_0[6]/m1_155_n223# dac_3v_cell_dummy_0[6]/m1_824_799#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[7] dac_3v_cell_dummy_0[7]/m4_99_18# dac_3v_cell_dummy_0[6]/w_316_892#
+ dac_3v_cell_dummy_0[7]/m4_99_276# dac_3v_cell_dummy_0[7]/m4_99_801# VSUBS dac_3v_cell_dummy_0[7]/m4_99_930#
+ dac_3v_cell_dummy_0[6]/m1_824_799# dac_3v_cell_dummy_0[7]/m4_99_405# dac_3v_cell_dummy_0[7]/m4_99_1059#
+ dac_3v_cell_dummy_0[7]/m4_99_672# dac_3v_cell_dummy_0[7]/w_316_892# dac_3v_cell_dummy_0[8]/m1_155_n223#
+ dac_3v_cell_dummy_0[7]/m4_99_147# dac_3v_cell_dummy_0[7]/m1_155_n223# dac_3v_cell_dummy_0[7]/m1_824_799#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[8] dac_3v_cell_dummy_0[8]/m4_99_18# dac_3v_cell_dummy_0[7]/w_316_892#
+ dac_3v_cell_dummy_0[8]/m4_99_276# dac_3v_cell_dummy_0[8]/m4_99_801# VSUBS dac_3v_cell_dummy_0[8]/m4_99_930#
+ dac_3v_cell_dummy_0[7]/m1_824_799# dac_3v_cell_dummy_0[8]/m4_99_405# dac_3v_cell_dummy_0[8]/m4_99_1059#
+ dac_3v_cell_dummy_0[8]/m4_99_672# dac_3v_cell_dummy_0[8]/w_316_892# m1_36_13186#
+ dac_3v_cell_dummy_0[8]/m4_99_147# dac_3v_cell_dummy_0[8]/m1_155_n223# m1_36_13186#
+ dac_3v_cell_dummy
Xdac_3v_cell_dummy_0[9] dac_3v_cell_dummy_0[9]/m4_99_18# dac_3v_cell_dummy_0[8]/w_316_892#
+ dac_3v_cell_dummy_0[9]/m4_99_276# dac_3v_cell_dummy_0[9]/m4_99_801# VSUBS dac_3v_cell_dummy_0[9]/m4_99_930#
+ m1_36_13186# dac_3v_cell_dummy_0[9]/m4_99_405# dac_3v_cell_dummy_0[9]/m4_99_1059#
+ dac_3v_cell_dummy_0[9]/m4_99_672# dac_3v_cell_dummy_0[9]/w_316_892# m1_28_15111#
+ dac_3v_cell_dummy_0[9]/m4_99_147# m1_36_13186# m1_28_15111# dac_3v_cell_dummy
.ends

.subckt sky130_ef_ip__rdac3v_8bit b0 b1 b2 b3 b4 b5 b6 b7 out vdd ena dvdd Vhigh Vlow
+ vss dvss
Xdac_3v_column_odd_0 b6b dac_3v_column_0/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a b6a b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a dac_3v_column_1/out_5 b1b b1b b3a vdd vdd
+ dac_3v_column_0/dum1_out b0a b1a dac_3v_column_1/res0_in b0b b2b b2a dac_3v_column_0/out_4
+ b1a vdd b2b b3b vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_2/in_5
+ b0a dac_3v_column_1/dum0_in b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xdac_3v_column_odd_1 b7b dac_3v_column_1/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a b7a b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a out_unbuf b1b b1b b3a vdd vdd dac_3v_column_1/dum1_out
+ b0a b1a dac_3v_column_2/res0_in b0b b2b b2a dac_3v_column_1/out_4 b1a vdd b2b b3b
+ vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_2/in_5
+ b0a dac_3v_column_2/dum0_in b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xdac_3v_column_odd_2 b6a dac_3v_column_2/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a b6b b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a dac_3v_column_3/out_5 b1b b1b b3a vdd vdd
+ dac_3v_column_2/dum1_out b0a b1a dac_3v_column_3/res0_in b0b b2b b2a dac_3v_column_2/out_4
+ b1a vdd b2b b3b vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_2/in_5
+ b0a dac_3v_column_3/dum0_in b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xdac_3v_column_odd_3 vdd dac_3v_column_3/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a vss b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a dac_3v_column_odd_3/in_5 b1b b1b b3a vdd
+ vdd dac_3v_column_3/dum1_out b0a b1a dac_3v_column_4/res0_in b0b b2b b2a dac_3v_column_3/out_4
+ b1a vdd b2b b3b vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_3/in_5
+ b0a dac_3v_column_4/dum0_in b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xdac_3v_column_odd_4 b6b dac_3v_column_4/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a b6a b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a dac_3v_column_5/out_5 b1b b1b b3a vdd vdd
+ dac_3v_column_4/dum1_out b0a b1a dac_3v_column_5/res0_in b0b b2b b2a dac_3v_column_4/out_4
+ b1a vdd b2b b3b vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_6/in_5
+ b0a dac_3v_column_5/dum0_in b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xfollower_amp_0 vdd out ena out_unbuf dvss vss follower_amp
Xdac_3v_column_odd_5 b7a dac_3v_column_5/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a b7b b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a out_unbuf b1b b1b b3a vdd vdd dac_3v_column_5/dum1_out
+ b0a b1a dac_3v_column_6/res0_in b0b b2b b2a dac_3v_column_5/out_4 b1a vdd b2b b3b
+ vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_6/in_5
+ b0a dac_3v_column_6/dum0_in b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xdac_3v_column_odd_6 b6a dac_3v_column_6/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a b6b b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a dac_3v_column_7/out_5 b1b b1b b3a vdd vdd
+ dac_3v_column_6/dum1_out b0a b1a dac_3v_column_7/res0_in b0b b2b b2a dac_3v_column_6/out_4
+ b1a vdd b2b b3b vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_6/in_5
+ b0a dac_3v_column_7/dum0_in b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xdac_3v_column_odd_7 vdd dac_3v_column_7/res1_out b3b b0b b0b b5b b0b b0b b2a b4a
+ b4b b0a b2b b0b b1b vdd vdd b1b b0b b5a b1b b0b b0a b0a vss b0a b1b b0a b3a b2a
+ b0a b0a b0b b0a vdd b0a b0a b0b b0b b0a dac_3v_column_odd_7/in_5 b1b b1b b3a vdd
+ vdd dac_3v_column_7/dum1_out b0a b1a Vlow b0b b2b b2a dac_3v_column_7/out_4 b1a
+ vdd b2b b3b vdd b1a b0b b2b b1a b1a b1a b0b b1b b1a b0a vdd vdd b0b dac_3v_column_odd_7/in_5
+ b0a dac_3v_column_odd_7/dum_out1 b1b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column_odd
Xdac_3v_column_0 b4b dac_3v_column_0/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_0/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_1/out_5 b0a
+ dac_3v_column_0/out_4 b5b b0a b1a b0b b3b b3a b1a vdd b2b Vhigh b2b vdd b1a b0b
+ b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a dac_3v_column_0/res1_out
+ b5a b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xdac_3v_column_1 b4b dac_3v_column_1/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_1/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_1/out_5 b0a
+ dac_3v_column_1/out_4 b5a b0a b1a b0b b3b b3a b1a vdd b2b dac_3v_column_1/res0_in
+ b2b vdd b1a b0b b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a
+ dac_3v_column_1/res1_out b5b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xdac_3v_column_2 b4b dac_3v_column_2/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_2/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_3/out_5 b0a
+ dac_3v_column_2/out_4 b5b b0a b1a b0b b3b b3a b1a vdd b2b dac_3v_column_2/res0_in
+ b2b vdd b1a b0b b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a
+ dac_3v_column_2/res1_out b5a b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xdac_3v_column_3 b4b dac_3v_column_3/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_3/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_3/out_5 b0a
+ dac_3v_column_3/out_4 b5a b0a b1a b0b b3b b3a b1a vdd b2b dac_3v_column_3/res0_in
+ b2b vdd b1a b0b b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a
+ dac_3v_column_3/res1_out b5b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xdac_3v_column_4 b4b dac_3v_column_4/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_4/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_5/out_5 b0a
+ dac_3v_column_4/out_4 b5b b0a b1a b0b b3b b3a b1a vdd b2b dac_3v_column_4/res0_in
+ b2b vdd b1a b0b b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a
+ dac_3v_column_4/res1_out b5a b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xdac_3v_column_5 b4b dac_3v_column_5/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_5/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_5/out_5 b0a
+ dac_3v_column_5/out_4 b5a b0a b1a b0b b3b b3a b1a vdd b2b dac_3v_column_5/res0_in
+ b2b vdd b1a b0b b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a
+ dac_3v_column_5/res1_out b5b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xdac_3v_column_6 b4b dac_3v_column_6/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_6/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_7/out_5 b0a
+ dac_3v_column_6/out_4 b5b b0a b1a b0b b3b b3a b1a vdd b2b dac_3v_column_6/res0_in
+ b2b vdd b1a b0b b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a
+ dac_3v_column_6/res1_out b5a b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xdac_3v_column_7 b4b dac_3v_column_7/dum1_out b0b b0b b2a b5b b0b b0b b2a b3a b4a
+ b0a b2a b0b vdd dac_3v_column_7/dum0_in vdd b0a b0b b5a b1b b0a b1b vdd b0a b1b
+ b1b b1b b3b b0b b0a b1b b0a b0b vdd b0a b0a b0a b0b b0a dac_3v_column_7/out_5 b0a
+ dac_3v_column_7/out_4 b5a b0a b1a b0b b3b b3a b1a vdd b2b dac_3v_column_7/res0_in
+ b2b vdd b1a b0b b0b b2b b1a b0b b1a b1b b2b vdd b1b b1a b0a vdd vdd b0b b0a b1a
+ dac_3v_column_7/res1_out b5b b0b vdd b1a b0a b0a b0b vdd b2a vss dac_3v_column
Xlevel_shifter_array_0 b2b b6b b2a b3 b7 b6a b3b dvdd b0 b3a b0a b4 b7a b4b b4a b1
+ b0b b5 b1b b7b b5a b5b b2 b1a dvss b6 vdd level_shifter_array
Xdac_3v_column_dummy_0 Vhigh b0a vdd b0b b1b b0a vdd b2a vss vss b4b b1b b2a b1b b1a
+ b2b b2a b1a b1b b1a b3b b3a b1b b1a b2a b2b b1a vdd b1b b5b vss vss b2b b1a vdd
+ b0a b0b b0a vdd b0b b0a b0b vss b1a b0a b4a vdd b0b vdd vss b0a b0b vss b1b b0a
+ dac_3v_column_0/dum0_in b0b b0b b0a vdd b0a b0b vdd b0a b0b vdd b2b b3a vdd b0b
+ b0a b0b b0a vdd vdd b0b vss vdd vdd b0a b1a vdd vdd vss vdd b0b m1_6304_841# vdd
+ b0a b0b b3b m1_6304_841# b5a b0a b1b b0b dac_3v_column_dummy
Xdac_3v_column_dummy_1 m1_25325_837# b0a vdd b0b b1b b0a vdd b2a vss vss b4b b1b b2a
+ b1b b1a b2b b2a b1a b1b b1a b3b b3a b1b b1a b2a b2b b1a vdd b1b b5b vss vss b2b
+ b1a vdd b0a b0b b0a vdd b0b b0a b0b vss b1a b0a b4a vdd b0b vdd vss b0a b0b vss
+ b1b b0a m1_25325_837# b0b b0b b0a vdd b0a b0b vdd b0a b0b vdd b2b b3a vdd b0b b0a
+ b0b b0a vdd vdd b0b vss vdd vdd b0a b1a vdd vdd vss vdd b0b Vlow vdd b0a b0b b3b
+ dac_3v_column_odd_7/dum_out1 b5a b0a b1b b0b dac_3v_column_dummy
.ends

.subckt simple_switch_array_32 vdda0 left_lp_opamp_p simplest_analog_switch_ena1v8_0[1|0]/on
+ comp_p left_lp_opamp_n simplest_analog_switch_ena1v8_0[1|4]/on comp_n simplest_analog_switch_ena1v8_0[0|4]/on
+ simplest_analog_switch_ena1v8_0[0|6]/on simplest_analog_switch_ena1v8_0[0|5]/on
+ dac1 simplest_analog_switch_ena1v8_0[1|6]/on dac0 amuxbusB amuxbusA simplest_analog_switch_ena1v8_1[0|0]/on
+ simplest_analog_switch_ena1v8_1[1|3]/on simplest_analog_switch_ena1v8_1[1|4]/on
+ analog0 right_hgbw_opamp_p simplest_analog_switch_ena1v8_0[0|8]/on simplest_analog_switch_ena1v8_0[1|9]/on
+ right_hgbw_opamp_n simplest_analog_switch_ena1v8_0[0|2]/on left_hgbw_opamp_p simplest_analog_switch_ena1v8_0[0|7]/on
+ simplest_analog_switch_ena1v8_1[1|2]/on simplest_analog_switch_ena1v8_0[1|2]/on
+ left_hgbw_opamp_n simplest_analog_switch_ena1v8_1[0|5]/on simplest_analog_switch_ena1v8_1[0|3]/on
+ simplest_analog_switch_ena1v8_0[1|7]/on simplest_analog_switch_ena1v8_0[1|8]/on
+ right_instramp_p simplest_analog_switch_ena1v8_0[0|9]/on simplest_analog_switch_ena1v8_0[0|3]/on
+ right_instramp_n simplest_analog_switch_ena1v8_0[1|5]/on simplest_analog_switch_ena1v8_1[1|5]/on
+ ulpcomp_p simplest_analog_switch_ena1v8_0[1|1]/on simplest_analog_switch_ena1v8_1[0|2]/on
+ ulpcomp_n simplest_analog_switch_ena1v8_1[0|1]/on simplest_analog_switch_ena1v8_1[0|4]/on
+ right_lp_opamp_p simplest_analog_switch_ena1v8_0[0|1]/on left_instramp_p adc1 simplest_analog_switch_ena1v8_0[0|0]/on
+ right_lp_opamp_n simplest_analog_switch_ena1v8_1[1|1]/on adc0 vccd0 simplest_analog_switch_ena1v8_0[1|3]/on
+ left_instramp_n simplest_analog_switch_ena1v8_1[1|0]/on vssa0 analog1 vssd0
Xsimplest_analog_switch_ena1v8_0[0|0] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[0|0]/on
+ analog1 vssd0 right_instramp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[1|0] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[1|0]/on
+ analog0 vssd0 right_instramp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[0|1] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[0|1]/on
+ analog1 vssd0 right_hgbw_opamp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[1|1] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[1|1]/on
+ analog0 vssd0 right_hgbw_opamp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[0|2] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[0|2]/on
+ analog1 vssd0 right_lp_opamp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[1|2] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[1|2]/on
+ analog0 vssd0 right_lp_opamp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[0|3] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[0|3]/on
+ analog1 vssd0 left_lp_opamp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[1|3] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[1|3]/on
+ analog0 vssd0 left_lp_opamp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[0|4] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[0|4]/on
+ analog1 vssd0 left_hgbw_opamp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[1|4] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[1|4]/on
+ analog0 vssd0 left_hgbw_opamp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[0|5] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[0|5]/on
+ analog1 vssd0 left_instramp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[1|5] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[1|5]/on
+ analog0 vssd0 left_instramp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[0|6] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[0|6]/on
+ analog1 vssd0 ulpcomp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[1|6] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[1|6]/on
+ analog0 vssd0 ulpcomp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[0|7] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[0|7]/on
+ analog1 vssd0 comp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[1|7] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[1|7]/on
+ analog0 vssd0 comp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[0|8] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[0|8]/on
+ analog1 vssd0 adc0 simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[1|8] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[1|8]/on
+ analog0 vssd0 adc1 simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[0|9] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[0|9]/on
+ analog1 vssd0 dac0 simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_0[1|9] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_0[1|9]/on
+ analog0 vssd0 dac1 simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[0|0] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[0|0]/on
+ amuxbusB vssd0 right_instramp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1|0] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[1|0]/on
+ amuxbusA vssd0 right_instramp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[0|1] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[0|1]/on
+ amuxbusB vssd0 right_hgbw_opamp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1|1] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[1|1]/on
+ amuxbusA vssd0 right_hgbw_opamp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[0|2] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[0|2]/on
+ amuxbusB vssd0 right_lp_opamp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1|2] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[1|2]/on
+ amuxbusA vssd0 right_lp_opamp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[0|3] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[0|3]/on
+ amuxbusB vssd0 left_lp_opamp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1|3] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[1|3]/on
+ amuxbusA vssd0 left_lp_opamp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[0|4] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[0|4]/on
+ amuxbusB vssd0 left_hgbw_opamp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1|4] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[1|4]/on
+ amuxbusA vssd0 left_hgbw_opamp_p simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[0|5] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[0|5]/on
+ amuxbusB vssd0 left_instramp_n simplest_analog_switch_ena1v8
Xsimplest_analog_switch_ena1v8_1[1|5] vdda0 vccd0 vssa0 simplest_analog_switch_ena1v8_1[1|5]/on
+ amuxbusA vssd0 left_instramp_p simplest_analog_switch_ena1v8
.ends

.subckt bias_generator_be4 dvdd dvss lsxo_src_50 en_user2_trim_n en_hsxo_trim_p en_hsxo_bias
+ en_brnout_bias en_lp2_bias en_lp1_trim_p en_lp1_bias en_lsxo_bias en_comp_trim_n
+ en_hsxo_trim_n en_snk_test hgbw1_src_100 instr2_src_100 comp_src_400 user_src_50
+ test_src_500 hsxo_src_100 idac_src_1000 en_idac_bias en_user2_bias en_user1_bias
+ en_user2_trim_p en_src_test en_comp_bias en_instr2_trim_p en_comp_trim_p en_ov_bias
+ en_instr1_bias en_hgbw2_trim_p en_instr1_trim_p en_instr2_bias en_hgbw1_bias en_lp2_trim_p
+ en_hgbw1_trim_p en_hgbw2_bias brnout_src_200 bandgap_snk_250 avdd bias_nstack_0[9]/nbias
+ lp1_src_100 bias_pstack_0[9]/pbias instr1_src_100 user_src_150 lp2_src_100 hgbw2_src_100
+ bias_pstack_0[9]/pcasc ov_src_600 avss
Xsky130_fd_sc_hvl__inv_2_16 sky130_fd_sc_hvl__inv_2_16/A dvss dvss avdd avdd bias_pstack_0[9]/enb
+ sky130_fd_sc_hvl__inv_2
Xbias_nstack_0[0] bias_nstack_0[9]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[0]/vcasc
+ bias_nstack
Xbias_nstack_0[1] bias_nstack_0[9]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[1]/vcasc
+ bias_nstack
Xbias_nstack_0[2] bias_nstack_0[9]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[2]/vcasc
+ bias_nstack
Xbias_nstack_0[3] bias_nstack_0[9]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[3]/vcasc
+ bias_nstack
Xbias_nstack_0[4] bias_nstack_0[9]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[4]/vcasc
+ bias_nstack
Xbias_nstack_0[5] bias_nstack_0[9]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[5]/vcasc
+ bias_nstack
Xbias_nstack_0[6] bias_nstack_0[9]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[6]/vcasc
+ bias_nstack
Xbias_nstack_0[7] bias_nstack_0[9]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[7]/vcasc
+ bias_nstack
Xbias_nstack_0[8] bias_nstack_0[9]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[8]/vcasc
+ bias_nstack
Xbias_nstack_0[9] bias_nstack_0[9]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[9]/vcasc
+ bias_nstack
Xbias_nstack_0[10] bias_nstack_0[9]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[10]/vcasc
+ bias_nstack
Xbias_nstack_0[11] bias_nstack_0[9]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[11]/vcasc
+ bias_nstack
Xbias_nstack_0[12] bias_nstack_0[9]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[12]/vcasc
+ bias_nstack
Xbias_nstack_0[13] bias_nstack_0[9]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[13]/vcasc
+ bias_nstack
Xbias_nstack_0[14] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[14]/vcasc bias_nstack
Xbias_nstack_0[15] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[15]/vcasc bias_nstack
Xbias_nstack_0[16] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[16]/vcasc bias_nstack
Xbias_nstack_0[17] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[17]/vcasc bias_nstack
Xbias_nstack_0[18] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[18]/vcasc bias_nstack
Xbias_nstack_0[19] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[19]/vcasc bias_nstack
Xbias_nstack_0[20] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[20]/vcasc bias_nstack
Xbias_nstack_0[21] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[21]/vcasc bias_nstack
Xbias_nstack_0[22] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[22]/vcasc bias_nstack
Xbias_nstack_0[23] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[23]/vcasc bias_nstack
Xbias_nstack_0[24] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[24]/vcasc bias_nstack
Xbias_nstack_0[25] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[25]/vcasc bias_nstack
Xbias_nstack_0[26] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[26]/vcasc bias_nstack
Xbias_nstack_0[27] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[27]/vcasc bias_nstack
Xbias_nstack_0[28] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[28]/vcasc bias_nstack
Xbias_nstack_0[29] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[29]/vcasc bias_nstack
Xbias_nstack_0[30] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[30]/vcasc bias_nstack
Xbias_nstack_0[31] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[31]/vcasc bias_nstack
Xbias_nstack_0[32] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[32]/vcasc bias_nstack
Xbias_nstack_0[33] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[33]/vcasc bias_nstack
Xbias_nstack_0[34] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[34]/vcasc bias_nstack
Xbias_nstack_0[35] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[35]/vcasc bias_nstack
Xbias_nstack_0[36] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[36]/vcasc bias_nstack
Xbias_nstack_0[37] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[37]/vcasc bias_nstack
Xbias_nstack_0[38] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[38]/vcasc bias_nstack
Xbias_nstack_0[39] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[39]/vcasc bias_nstack
Xbias_nstack_0[40] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[40]/vcasc bias_nstack
Xbias_nstack_0[41] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[41]/vcasc bias_nstack
Xbias_nstack_0[42] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[42]/vcasc bias_nstack
Xbias_nstack_0[43] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[43]/vcasc bias_nstack
Xbias_nstack_0[44] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[44]/vcasc bias_nstack
Xbias_nstack_0[45] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[45]/vcasc bias_nstack
Xbias_nstack_0[46] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[46]/vcasc bias_nstack
Xbias_nstack_0[47] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[47]/vcasc bias_nstack
Xbias_nstack_0[48] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[48]/vcasc bias_nstack
Xbias_nstack_0[49] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[49]/vcasc bias_nstack
Xbias_nstack_0[50] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[50]/vcasc bias_nstack
Xbias_nstack_0[51] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[51]/vcasc bias_nstack
Xbias_nstack_0[52] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[52]/vcasc bias_nstack
Xbias_nstack_0[53] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[53]/vcasc bias_nstack
Xbias_nstack_0[54] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[54]/vcasc bias_nstack
Xbias_nstack_0[55] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[55]/vcasc bias_nstack
Xbias_nstack_0[56] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[56]/vcasc bias_nstack
Xbias_nstack_0[57] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[57]/vcasc bias_nstack
Xbias_nstack_0[58] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[58]/vcasc bias_nstack
Xbias_nstack_0[59] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[59]/vcasc bias_nstack
Xbias_nstack_0[60] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[60]/vcasc bias_nstack
Xbias_nstack_0[61] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[61]/vcasc bias_nstack
Xbias_nstack_0[62] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[62]/vcasc bias_nstack
Xbias_nstack_0[63] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[63]/vcasc bias_nstack
Xbias_nstack_0[64] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[64]/vcasc bias_nstack
Xbias_nstack_0[65] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[65]/vcasc bias_nstack
Xbias_nstack_0[66] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[66]/vcasc bias_nstack
Xbias_nstack_0[67] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[67]/vcasc bias_nstack
Xbias_nstack_0[68] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[68]/vcasc bias_nstack
Xbias_nstack_0[69] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[69]/vcasc bias_nstack
Xbias_nstack_0[70] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[70]/vcasc bias_nstack
Xbias_nstack_0[71] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[71]/vcasc bias_nstack
Xbias_nstack_0[72] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[72]/vcasc bias_nstack
Xbias_nstack_0[73] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[73]/vcasc bias_nstack
Xbias_nstack_0[74] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[74]/vcasc bias_nstack
Xbias_nstack_0[75] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[75]/vcasc bias_nstack
Xbias_nstack_0[76] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[76]/vcasc bias_nstack
Xbias_nstack_0[77] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[77]/vcasc bias_nstack
Xbias_nstack_0[78] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[78]/vcasc bias_nstack
Xbias_nstack_0[79] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[79]/vcasc bias_nstack
Xbias_nstack_0[80] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[80]/vcasc bias_nstack
Xbias_nstack_0[81] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[81]/vcasc bias_nstack
Xbias_nstack_0[82] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[82]/vcasc bias_nstack
Xbias_nstack_0[83] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[83]/vcasc bias_nstack
Xbias_nstack_0[84] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[84]/vcasc bias_nstack
Xbias_nstack_0[85] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[85]/vcasc bias_nstack
Xbias_nstack_0[86] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[86]/vcasc bias_nstack
Xbias_nstack_0[87] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[87]/vcasc bias_nstack
Xbias_nstack_0[88] test_src_500 bias_nstack_0[88]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[88]/vcasc bias_nstack
Xbias_nstack_0[89] bandgap_snk_250 bias_nstack_0[93]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[89]/vcasc bias_nstack
Xbias_nstack_0[90] bandgap_snk_250 bias_nstack_0[93]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[90]/vcasc bias_nstack
Xbias_nstack_0[91] bandgap_snk_250 bias_nstack_0[93]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[91]/vcasc bias_nstack
Xbias_nstack_0[92] bandgap_snk_250 bias_nstack_0[93]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[92]/vcasc bias_nstack
Xbias_nstack_0[93] bandgap_snk_250 bias_nstack_0[93]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[93]/vcasc bias_nstack
Xbias_nstack_0[94] user_src_150 bias_nstack_0[95]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[94]/vcasc bias_nstack
Xbias_nstack_0[95] user_src_150 bias_nstack_0[95]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[95]/vcasc bias_nstack
Xbias_nstack_0[96] comp_src_400 bias_nstack_0[97]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[96]/vcasc bias_nstack
Xbias_nstack_0[97] comp_src_400 bias_nstack_0[97]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[97]/vcasc bias_nstack
Xbias_nstack_0[98] hsxo_src_100 bias_nstack_0[99]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[98]/vcasc bias_nstack
Xbias_nstack_0[99] hsxo_src_100 bias_nstack_0[99]/ena bias_nstack_0[9]/nbias avss
+ bias_nstack_0[99]/vcasc bias_nstack
Xbias_nstack_0[100] bias_nstack_0[101]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[100]/vcasc
+ bias_nstack
Xbias_nstack_0[101] bias_nstack_0[101]/itail avss bias_nstack_0[9]/nbias avss bias_nstack_0[101]/vcasc
+ bias_nstack
Xsky130_fd_sc_hvl__inv_2_17 sky130_fd_sc_hvl__inv_2_17/A dvss dvss avdd avdd bias_pstack_0[40]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_18 sky130_fd_sc_hvl__inv_2_18/A dvss dvss avdd avdd bias_pstack_0[44]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_19 sky130_fd_sc_hvl__inv_2_19/A dvss dvss avdd avdd bias_pstack_0[38]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_0 sky130_fd_sc_hvl__inv_2_0/A dvss dvss avdd avdd bias_pstack_0[95]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_1 sky130_fd_sc_hvl__inv_2_1/A dvss dvss avdd avdd bias_pstack_0[90]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_20 en_comp_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_2_2 sky130_fd_sc_hvl__inv_2_2/A dvss dvss avdd avdd bias_pstack_0[80]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_10 en_lp1_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_21 en_instr1_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|0] en_snk_test dvdd dvss avdd avdd bias_nstack_0[88]/ena
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|0] en_user2_trim_n dvdd dvss avdd avdd bias_nstack_0[95]/ena
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[2|0] en_comp_trim_n dvdd dvss avdd avdd bias_nstack_0[97]/ena
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[3|0] en_hsxo_trim_n dvdd dvss avdd avdd bias_nstack_0[99]/ena
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|1] en_lp2_bias dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_0/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|1] en_lp1_trim_p dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_7/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[2|1] en_lsxo_bias dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_11/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[3|1] en_lp1_bias dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_10/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|2] en_hgbw2_bias dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_12/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|2] en_hgbw1_trim_p dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_1/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[2|2] en_lp2_trim_p dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_6/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[3|2] en_hgbw1_bias dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_5/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|3] en_instr2_bias dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_8/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|3] en_instr1_trim_p dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_13/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[2|3] en_hgbw2_trim_p dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_14/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[3|3] en_instr1_bias dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_15/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|4] en_ov_bias dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_9/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|4] en_comp_trim_p dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_4/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[2|4] en_instr2_trim_p dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_3/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[3|4] en_comp_bias dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_2/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|5] en_src_test dvdd dvss avdd avdd bias_nstack_0[93]/ena
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|5] en_user2_trim_p dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_23/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[2|5] en_user1_bias dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_22/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[3|5] en_user2_bias dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_21/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[0|6] en_idac_bias dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_16/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[1|6] en_hsxo_trim_p dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_19/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[2|6] en_brnout_bias dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_18/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__lsbuflv2hv_1_0[3|6] en_hsxo_bias dvdd dvss avdd avdd sky130_fd_sc_hvl__inv_2_17/A
+ avdd dvss dvss sky130_fd_sc_hvl__lsbuflv2hv_1
Xsky130_fd_sc_hvl__inv_2_3 sky130_fd_sc_hvl__inv_2_3/A dvss dvss avdd avdd bias_pstack_0[81]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_11 en_hgbw1_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_22 en_hgbw1_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_2_4 sky130_fd_sc_hvl__inv_2_4/A dvss dvss avdd avdd bias_pstack_0[72]/enb
+ sky130_fd_sc_hvl__inv_2
Xbias_pstack_0[0] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[0]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[1] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[1]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[2] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[2]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[3] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[3]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[4] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[4]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[5] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[5]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[6] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[6]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[7] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[7]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[8] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[8]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[9] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[9]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[10] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[10]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[11] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[11]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[12] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[12]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[13] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[13]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[14] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[14]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[15] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[15]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[16] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[16]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[17] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[17]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[18] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[18]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[19] bias_pstack_0[9]/pcasc bias_pstack_0[9]/enb idac_src_1000 bias_pstack_0[19]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[20] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[20]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[21] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[21]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[22] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[22]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[23] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[23]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[24] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[24]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[25] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[25]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[26] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[26]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[27] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[27]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[28] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[28]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[29] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[29]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[30] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[30]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[31] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[31]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[32] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[32]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[33] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[33]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[34] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[34]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[35] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[35]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[36] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[36]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[37] bias_pstack_0[9]/pcasc avdd bias_pstack_0[37]/itail bias_pstack_0[37]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[38] bias_pstack_0[9]/pcasc bias_pstack_0[38]/enb hsxo_src_100 bias_pstack_0[38]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[39] bias_pstack_0[9]/pcasc bias_pstack_0[40]/enb hsxo_src_100 bias_pstack_0[39]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[40] bias_pstack_0[9]/pcasc bias_pstack_0[40]/enb hsxo_src_100 bias_pstack_0[40]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[41] bias_pstack_0[9]/pcasc bias_pstack_0[44]/enb brnout_src_200 bias_pstack_0[41]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[42] bias_pstack_0[9]/pcasc bias_pstack_0[44]/enb brnout_src_200 bias_pstack_0[42]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[43] bias_pstack_0[9]/pcasc bias_pstack_0[44]/enb brnout_src_200 bias_pstack_0[43]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[44] bias_pstack_0[9]/pcasc bias_pstack_0[44]/enb brnout_src_200 bias_pstack_0[44]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[45] bias_pstack_0[9]/pcasc bias_pstack_0[54]/enb test_src_500 bias_pstack_0[45]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[46] bias_pstack_0[9]/pcasc bias_pstack_0[54]/enb test_src_500 bias_pstack_0[46]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[47] bias_pstack_0[9]/pcasc bias_pstack_0[54]/enb test_src_500 bias_pstack_0[47]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[48] bias_pstack_0[9]/pcasc bias_pstack_0[54]/enb test_src_500 bias_pstack_0[48]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[49] bias_pstack_0[9]/pcasc bias_pstack_0[54]/enb test_src_500 bias_pstack_0[49]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[50] bias_pstack_0[9]/pcasc bias_pstack_0[54]/enb test_src_500 bias_pstack_0[50]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[51] bias_pstack_0[9]/pcasc bias_pstack_0[54]/enb test_src_500 bias_pstack_0[51]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[52] bias_pstack_0[9]/pcasc bias_pstack_0[54]/enb test_src_500 bias_pstack_0[52]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[53] bias_pstack_0[9]/pcasc bias_pstack_0[54]/enb test_src_500 bias_pstack_0[53]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[54] bias_pstack_0[9]/pcasc bias_pstack_0[54]/enb test_src_500 bias_pstack_0[54]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[55] bias_pstack_0[9]/pcasc bias_pstack_0[55]/enb user_src_150 bias_pstack_0[55]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[56] bias_pstack_0[9]/pcasc bias_pstack_0[58]/enb user_src_150 bias_pstack_0[56]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[57] bias_pstack_0[9]/pcasc bias_pstack_0[58]/enb user_src_150 bias_pstack_0[57]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[58] bias_pstack_0[9]/pcasc bias_pstack_0[58]/enb user_src_150 bias_pstack_0[58]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[59] bias_pstack_0[9]/pcasc bias_pstack_0[59]/enb user_src_50 bias_pstack_0[59]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[60] bias_pstack_0[9]/pcasc bias_pstack_0[71]/enb ov_src_600 bias_pstack_0[60]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[61] bias_pstack_0[9]/pcasc bias_pstack_0[71]/enb ov_src_600 bias_pstack_0[61]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[62] bias_pstack_0[9]/pcasc bias_pstack_0[71]/enb ov_src_600 bias_pstack_0[62]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[63] bias_pstack_0[9]/pcasc bias_pstack_0[71]/enb ov_src_600 bias_pstack_0[63]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[64] bias_pstack_0[9]/pcasc bias_pstack_0[71]/enb ov_src_600 bias_pstack_0[64]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[65] bias_pstack_0[9]/pcasc bias_pstack_0[71]/enb ov_src_600 bias_pstack_0[65]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[66] bias_pstack_0[9]/pcasc bias_pstack_0[71]/enb ov_src_600 bias_pstack_0[66]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[67] bias_pstack_0[9]/pcasc bias_pstack_0[71]/enb ov_src_600 bias_pstack_0[67]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[68] bias_pstack_0[9]/pcasc bias_pstack_0[71]/enb ov_src_600 bias_pstack_0[68]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[69] bias_pstack_0[9]/pcasc bias_pstack_0[71]/enb ov_src_600 bias_pstack_0[69]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[70] bias_pstack_0[9]/pcasc bias_pstack_0[71]/enb ov_src_600 bias_pstack_0[70]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[71] bias_pstack_0[9]/pcasc bias_pstack_0[71]/enb ov_src_600 bias_pstack_0[71]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[72] bias_pstack_0[9]/pcasc bias_pstack_0[72]/enb comp_src_400 bias_pstack_0[72]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[73] bias_pstack_0[9]/pcasc bias_pstack_0[80]/enb comp_src_400 bias_pstack_0[73]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[74] bias_pstack_0[9]/pcasc bias_pstack_0[80]/enb comp_src_400 bias_pstack_0[74]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[75] bias_pstack_0[9]/pcasc bias_pstack_0[80]/enb comp_src_400 bias_pstack_0[75]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[76] bias_pstack_0[9]/pcasc bias_pstack_0[80]/enb comp_src_400 bias_pstack_0[76]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[77] bias_pstack_0[9]/pcasc bias_pstack_0[80]/enb comp_src_400 bias_pstack_0[77]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[78] bias_pstack_0[9]/pcasc bias_pstack_0[80]/enb comp_src_400 bias_pstack_0[78]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[79] bias_pstack_0[9]/pcasc bias_pstack_0[80]/enb comp_src_400 bias_pstack_0[79]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[80] bias_pstack_0[9]/pcasc bias_pstack_0[80]/enb comp_src_400 bias_pstack_0[80]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[81] bias_pstack_0[9]/pcasc bias_pstack_0[81]/enb instr2_src_100 bias_pstack_0[81]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[82] bias_pstack_0[9]/pcasc bias_pstack_0[83]/enb instr2_src_100 bias_pstack_0[82]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[83] bias_pstack_0[9]/pcasc bias_pstack_0[83]/enb instr2_src_100 bias_pstack_0[83]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[84] bias_pstack_0[9]/pcasc bias_pstack_0[84]/enb instr1_src_100 bias_pstack_0[84]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[85] bias_pstack_0[9]/pcasc bias_pstack_0[86]/enb instr1_src_100 bias_pstack_0[85]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[86] bias_pstack_0[9]/pcasc bias_pstack_0[86]/enb instr1_src_100 bias_pstack_0[86]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[87] bias_pstack_0[9]/pcasc bias_pstack_0[87]/enb hgbw2_src_100 bias_pstack_0[87]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[88] bias_pstack_0[9]/pcasc bias_pstack_0[89]/enb hgbw2_src_100 bias_pstack_0[88]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[89] bias_pstack_0[9]/pcasc bias_pstack_0[89]/enb hgbw2_src_100 bias_pstack_0[89]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[90] bias_pstack_0[9]/pcasc bias_pstack_0[90]/enb hgbw1_src_100 bias_pstack_0[90]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[91] bias_pstack_0[9]/pcasc bias_pstack_0[92]/enb hgbw1_src_100 bias_pstack_0[91]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[92] bias_pstack_0[9]/pcasc bias_pstack_0[92]/enb hgbw1_src_100 bias_pstack_0[92]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[93] bias_pstack_0[9]/pcasc bias_pstack_0[93]/enb lp2_src_100 bias_pstack_0[93]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[94] bias_pstack_0[9]/pcasc bias_pstack_0[95]/enb lp2_src_100 bias_pstack_0[94]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[95] bias_pstack_0[9]/pcasc bias_pstack_0[95]/enb lp2_src_100 bias_pstack_0[95]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[96] bias_pstack_0[9]/pcasc bias_pstack_0[96]/enb lp1_src_100 bias_pstack_0[96]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[97] bias_pstack_0[9]/pcasc bias_pstack_0[98]/enb lp1_src_100 bias_pstack_0[97]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[98] bias_pstack_0[9]/pcasc bias_pstack_0[98]/enb lp1_src_100 bias_pstack_0[98]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[99] bias_pstack_0[9]/pcasc bias_pstack_0[99]/enb lsxo_src_50 bias_pstack_0[99]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[100] bias_pstack_0[9]/pcasc avdd bias_pstack_0[101]/itail bias_pstack_0[100]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xbias_pstack_0[101] bias_pstack_0[9]/pcasc avdd bias_pstack_0[101]/itail bias_pstack_0[101]/vcasc
+ bias_pstack_0[9]/pbias avss avdd bias_pstack
Xsky130_fd_sc_hvl__diode_2_12 en_instr1_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_23 en_lp1_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_2_5 sky130_fd_sc_hvl__inv_2_5/A dvss dvss avdd avdd bias_pstack_0[92]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_13 en_comp_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_24 en_lp2_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_2_6 sky130_fd_sc_hvl__inv_2_6/A dvss dvss avdd avdd bias_pstack_0[93]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_14 en_user2_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_25 en_hgbw2_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_2_7 sky130_fd_sc_hvl__inv_2_7/A dvss dvss avdd avdd bias_pstack_0[96]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_15 en_lsxo_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_26 en_instr2_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_2_8 sky130_fd_sc_hvl__inv_2_8/A dvss dvss avdd avdd bias_pstack_0[83]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_16 en_hsxo_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_27 en_user1_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_2_9 sky130_fd_sc_hvl__inv_2_9/A dvss dvss avdd avdd bias_pstack_0[71]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_17 en_brnout_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_18 en_hsxo_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_19 en_user2_trim_p dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_0 en_snk_test dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_1 en_idac_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_2 en_src_test dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_14 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_3 en_ov_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_4 en_instr2_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__diode_2_5 en_hgbw2_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_2_20 bias_nstack_0[93]/ena dvss dvss avdd avdd bias_pstack_0[54]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_6 en_lp2_bias dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_18 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__inv_2_21 sky130_fd_sc_hvl__inv_2_21/A dvss dvss avdd avdd bias_pstack_0[58]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_10 sky130_fd_sc_hvl__inv_2_10/A dvss dvss avdd avdd bias_pstack_0[98]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__decap_4_0 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__diode_2_7 en_comp_trim_n dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__decap_4_1 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
Xsky130_fd_sc_hvl__inv_2_22 sky130_fd_sc_hvl__inv_2_22/A dvss dvss avdd avdd bias_pstack_0[59]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_11 sky130_fd_sc_hvl__inv_2_11/A dvss dvss avdd avdd bias_pstack_0[99]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_8 en_user2_trim_n dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_2_23 sky130_fd_sc_hvl__inv_2_23/A dvss dvss avdd avdd bias_pstack_0[55]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_12 sky130_fd_sc_hvl__inv_2_12/A dvss dvss avdd avdd bias_pstack_0[89]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__diode_2_9 en_hsxo_trim_n dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
Xsky130_fd_sc_hvl__inv_2_13 sky130_fd_sc_hvl__inv_2_13/A dvss dvss avdd avdd bias_pstack_0[84]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_14 sky130_fd_sc_hvl__inv_2_14/A dvss dvss avdd avdd bias_pstack_0[87]/enb
+ sky130_fd_sc_hvl__inv_2
Xsky130_fd_sc_hvl__inv_2_15 sky130_fd_sc_hvl__inv_2_15/A dvss dvss avdd avdd bias_pstack_0[86]/enb
+ sky130_fd_sc_hvl__inv_2
.ends

.subckt sky130_ef_ip__biasgen4 ena ref_sel_vbg dvdd avdd vbg en_snk_test en_user2_trim_n
+ en_comp_trim_n en_hsxo_trim_n en_lp2_bias en_lp1_trim_p en_lsxo_bias en_lp1_bias
+ en_hgbw1_trim_p en_lp2_trim_p en_hgbw1_bias en_instr2_bias en_instr1_trim_p en_hgbw2_trim_p
+ en_instr1_bias en_ov_bias en_comp_trim_p en_instr2_trim_p en_comp_bias en_src_test
+ en_user2_trim_p en_user1_bias en_user2_bias en_idac_bias en_hsxo_trim_p en_brnout_bias
+ en_hsxo_bias en_hgbw2_bias lsxo_src_50 lp1_src_100 lp2_src_100 hgbw1_src_100 hgbw2_src_100
+ instr1_src_100 instr2_src_100 ov_src_600 user_src_50 test_src_500 brnout_src_200
+ hsxo_src_100 idac_src_1000 ref_in comp_src_400 bandgap_snk_250 user_src_150 dvss
+ avss
Xbias_generator_be4_0 dvdd dvss lsxo_src_50 en_user2_trim_n en_hsxo_trim_p en_hsxo_bias
+ en_brnout_bias en_lp2_bias en_lp1_trim_p en_lp1_bias en_lsxo_bias en_comp_trim_n
+ en_hsxo_trim_n en_snk_test hgbw1_src_100 instr2_src_100 comp_src_400 user_src_50
+ test_src_500 hsxo_src_100 idac_src_1000 en_idac_bias en_user2_bias en_user1_bias
+ en_user2_trim_p en_src_test en_comp_bias en_instr2_trim_p en_comp_trim_p en_ov_bias
+ en_instr1_bias en_hgbw2_trim_p en_instr1_trim_p en_instr2_bias en_hgbw1_bias en_lp2_trim_p
+ en_hgbw1_trim_p en_hgbw2_bias brnout_src_200 bandgap_snk_250 avdd bias_generator_fe_0/bias_amp_0/nbias
+ lp1_src_100 bias_generator_fe_0/bias_amp_0/out instr1_src_100 user_src_150 lp2_src_100
+ hgbw2_src_100 bias_generator_fe_0/bias_pstack_0[9]/pcasc ov_src_600 avss bias_generator_be4
Xbias_generator_fe_0 bias_generator_fe_0/snk_test0 bias_generator_fe_0/src_test0 vbg
+ ref_in dvss dvss ref_sel_vbg dvdd dvss bias_generator_fe_0/bias_amp_0/out avdd bias_generator_fe_0/bias_amp_0/nbias
+ ena bias_generator_fe_0/bias_pstack_0[9]/pcasc avss bias_generator_fe
.ends

.subckt bg__cap c1_n1050_n1000# m3_n1150_n1100#
X0 c1_n1050_n1000# m3_n1150_n1100# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
.ends

.subckt bg__res a_n1613_1296# a_n455_n1732# a_n3157_n1732# a_1089_n1732# a_n1227_n1732#
+ a_317_1296# a_n2771_n1732# a_703_1296# a_2247_n1732# a_2247_1296# a_2633_1296# a_n69_n1732#
+ a_n3929_n1732# a_3791_n1732# a_n2385_1296# a_1861_n1732# a_703_n1732# a_n2771_1296#
+ a_n3929_1296# a_3405_n1732# a_n69_1296# a_n455_1296# a_n841_1296# a_n2385_n1732#
+ a_n1999_1296# a_n1999_n1732# a_3019_1296# a_3405_1296# a_n841_n1732# a_n3543_n1732#
+ a_3791_1296# a_1475_n1732# a_317_n1732# a_n1613_n1732# a_n3157_1296# a_3019_n1732#
+ a_1089_1296# a_n3543_1296# a_1475_1296# a_2633_n1732# a_1861_1296# a_n4059_n1862#
+ a_n1227_1296#
X0 a_317_1296# a_317_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X1 a_n69_1296# a_n69_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X2 a_1861_1296# a_1861_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X3 a_703_1296# a_703_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X4 a_n2385_1296# a_n2385_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X5 a_n1227_1296# a_n1227_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X6 a_2247_1296# a_2247_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X7 a_n1999_1296# a_n1999_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X8 a_n1613_1296# a_n1613_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X9 a_n2771_1296# a_n2771_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X10 a_2633_1296# a_2633_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X11 a_3791_1296# a_3791_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X12 a_n3157_1296# a_n3157_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X13 a_3019_1296# a_3019_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X14 a_n3543_1296# a_n3543_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X15 a_3405_1296# a_3405_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X16 a_n455_1296# a_n455_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X17 a_1089_1296# a_1089_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X18 a_n841_1296# a_n841_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X19 a_n3929_1296# a_n3929_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
X20 a_1475_1296# a_1475_n1732# a_n4059_n1862# sky130_fd_pr__res_xhigh_po_0p69 l=13.12
.ends

.subckt bgt__MN a_n108_n231# a_n210_n343# a_50_n231# a_n50_n257#
X0 a_50_n231# a_n50_n257# a_n108_n231# a_n210_n343# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
.ends

.subckt bgt__res a_n1996_n712# a_n3056_n712# a_124_276# a_n936_276# a_1714_276# a_1714_n712#
+ a_n2526_276# a_654_276# a_n1466_n712# a_n1466_276# a_n4116_n712# a_n4246_n842# a_3304_276#
+ a_2244_276# a_1184_n712# a_n4116_276# a_2774_n712# a_1184_276# a_n3056_276# a_n1996_276#
+ a_3834_276# a_n2526_n712# a_2774_276# a_654_n712# a_3834_n712# a_2244_n712# a_n936_n712#
+ a_n3586_276# a_n3586_n712# a_n406_276# a_124_n712# a_n406_n712# a_3304_n712#
X0 a_n3586_276# a_n3586_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X1 a_n1466_276# a_n1466_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X2 a_3834_276# a_3834_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X3 a_1714_276# a_1714_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X4 a_n936_276# a_n936_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X5 a_n3056_276# a_n3056_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X6 a_2774_276# a_2774_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X7 a_3304_276# a_3304_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X8 a_n406_276# a_n406_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X9 a_2244_276# a_2244_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X10 a_1184_276# a_1184_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X11 a_654_276# a_654_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X12 a_124_276# a_124_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X13 a_n2526_276# a_n2526_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X14 a_n1996_276# a_n1996_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
X15 a_n4116_276# a_n4116_n712# a_n4246_n842# sky130_fd_pr__res_high_po_1p41 l=2.92
.ends

.subckt bg__trim m2_4223_3828# m2_800_5948# m2_640_4888# m2_4223_648# bgt__res_0/a_3834_n712#
+ m2_1120_8068# m2_480_3828# m2_4223_2768# m2_320_2768# m1_4339_1060# m1_1336_1060#
+ m2_4223_5948# m2_4223_8068# m2_160_1708# m1_3744_8480# m2_4223_4888# m2_4223_1708#
+ m2_960_7008# m2_0_648# VSUBS m2_4223_7008#
Xbgt__MN_0 m1_4339_1060# VSUBS m1_3744_8480# m2_4223_8068# bgt__MN
Xbgt__MN_1 m1_4339_1060# VSUBS m1_3323_1060# m2_4223_648# bgt__MN
Xbgt__MN_2 m1_4339_1060# VSUBS m1_3323_2120# m2_4223_1708# bgt__MN
Xbgt__MN_3 m1_4339_1060# VSUBS m1_3323_3180# m2_4223_2768# bgt__MN
Xbgt__MN_5 m1_4339_1060# VSUBS m1_3323_5300# m2_4223_4888# bgt__MN
Xbgt__MN_4 m1_4339_1060# VSUBS m1_3323_4240# m2_4223_3828# bgt__MN
Xbgt__MN_6 m1_1336_1060# VSUBS m1_1849_8480# m2_1120_8068# bgt__MN
Xbgt__MN_7 m1_4339_1060# VSUBS m1_3323_6360# m2_4223_5948# bgt__MN
Xbgt__MN_8 m1_4339_1060# VSUBS m1_3323_7420# m2_4223_7008# bgt__MN
Xbgt__MN_9 m1_1336_1060# VSUBS m1_1849_1060# m2_0_648# bgt__MN
Xbgt__MN_10 m1_1336_1060# VSUBS m1_1849_2120# m2_160_1708# bgt__MN
Xbgt__MN_11 m1_1336_1060# VSUBS m1_1849_3180# m2_320_2768# bgt__MN
Xbgt__MN_12 m1_1336_1060# VSUBS m1_1849_4240# m2_480_3828# bgt__MN
Xbgt__MN_13 m1_1336_1060# VSUBS m1_1849_5300# m2_640_4888# bgt__MN
Xbgt__MN_14 m1_1336_1060# VSUBS m1_1849_6360# m2_800_5948# bgt__MN
Xbgt__MN_15 m1_1336_1060# VSUBS m1_1849_7420# m2_960_7008# bgt__MN
Xbgt__res_0 m1_3323_6360# m1_3323_7420# m1_1849_4240# m1_1849_5300# m1_1849_3180#
+ m1_3323_2120# m1_1849_7420# m1_1849_4240# m1_3323_5300# m1_1849_6360# m1_3744_8480#
+ VSUBS m1_1849_1060# m1_1849_2120# m1_3323_3180# m1_1849_8480# m1_3323_1060# m1_1849_3180#
+ m1_1849_7420# m1_1849_6360# m1_1849_1060# m1_3323_6360# m1_1849_2120# m1_3323_3180#
+ bgt__res_0/a_3834_n712# m1_3323_2120# m1_3323_5300# m1_1849_8480# m1_3323_7420#
+ m1_1849_5300# m1_3323_4240# m1_3323_4240# m1_3323_1060# bgt__res
.ends

.subckt bgs__M3_M4 a_n287_n131# a_29_n157# a_229_n131# a_n229_n157# a_n389_n243# a_n29_n131#
X0 a_n29_n131# a_n229_n157# a_n287_n131# a_n389_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1 a_229_n131# a_29_n157# a_n29_n131# a_n389_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
.ends

.subckt bgs__M5_M6 w_n425_n284# a_n287_n136# a_229_n136# a_29_n162# a_n29_n136# a_n229_n162#
X0 a_n29_n136# a_n229_n162# a_n287_n136# w_n425_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X1 a_229_n136# a_29_n162# a_n29_n136# w_n425_n284# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
.ends

.subckt bgs__M7 a_100_n136# w_n296_n284# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n296_n284# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bg__startup m2_545_805# VSUBS m1_453_173# bgs__M5_M6_0/w_n425_n284# m2_1443_341#
+ m1_3178_549# m1_1258_542# bgs__M7_0/w_n296_n284# bgs__M3_M4_0/a_n287_n131# bgs__M7_0/a_100_n136#
Xbgs__M3_M4_0 bgs__M3_M4_0/a_n287_n131# m2_545_805# m1_251_542# m1_251_542# VSUBS
+ m1_453_173# bgs__M3_M4
Xbgs__M5_M6_0 bgs__M5_M6_0/w_n425_n284# m1_251_542# m1_1258_542# m1_1258_542# m2_1443_341#
+ m1_1258_542# bgs__M5_M6
Xbgs__M7_0 bgs__M7_0/a_100_n136# bgs__M7_0/w_n296_n284# m1_1258_542# m1_3178_549#
+ bgs__M7
.ends

.subckt bg__M1_M2 a_n287_n436# a_n487_n462# w_n683_n584# a_229_n436# a_29_n462# a_n545_n436#
+ a_n29_n436# a_n229_n462# a_487_n436# a_287_n462#
X0 a_n287_n436# a_n487_n462# a_n545_n436# w_n683_n584# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X1 a_487_n436# a_287_n462# a_229_n436# w_n683_n584# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X2 a_229_n436# a_29_n462# a_n29_n436# w_n683_n584# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 a_n29_n436# a_n229_n462# a_n287_n436# w_n683_n584# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
.ends

.subckt bgpg__pnp a_26_26# w_153_153# a_330_330#
X0 a_26_26# w_153_153# a_330_330# sky130_fd_pr__pnp_05v5_W0p68L0p68
**devattr s=18496,544
.ends

.subckt bg__pnp_group eg eu VDD GND
Xbgpg__pnp_0 GND GND eg bgpg__pnp
Xbgpg__pnp_1 GND GND eg bgpg__pnp
Xbgpg__pnp_2 GND GND eg bgpg__pnp
Xbgpg__pnp_3 GND GND eg bgpg__pnp
Xbgpg__pnp_4 GND GND eg bgpg__pnp
Xbgpg__pnp_5 GND GND eg bgpg__pnp
Xbgpg__pnp_6 GND GND eu bgpg__pnp
Xbgpg__pnp_7 GND GND eg bgpg__pnp
Xbgpg__pnp_8 GND GND eg bgpg__pnp
.ends

.subckt bgfcpm__DUM w_n194_n198# a_100_n136# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n194_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfcpm__M1 w_n194_n198# a_100_n136# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n194_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfcpm__MB2 w_n194_n198# a_100_n136# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n194_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfcpm__MB3 w_n194_n198# a_100_n136# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n194_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfc__pmirr vbp1 diff vbn2 vdd
Xbgfcpm__DUM_3 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_28 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_17 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_4 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__M1_0 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__DUM_29 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_18 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_5 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__M1_1 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__DUM_19 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_6 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__M1_2 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__DUM_7 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__M1_3 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__M1_4 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__DUM_8 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__M1_5 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__DUM_9 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__M1_6 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__M1_7 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__M1_8 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__M1_9 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__MB2_0 vdd vdd vbp1 vbp1 bgfcpm__MB2
Xbgfcpm__M1_10 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__MB2_1 vdd vdd vbp1 vbp1 bgfcpm__MB2
Xbgfcpm__M1_11 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__MB2_2 vdd vbp1 vdd vbp1 bgfcpm__MB2
Xbgfcpm__M1_12 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__MB2_3 vdd vbp1 vdd vbp1 bgfcpm__MB2
Xbgfcpm__M1_13 vdd vdd diff vbp1 bgfcpm__M1
Xbgfcpm__M1_14 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__M1_15 vdd diff vdd vbp1 bgfcpm__M1
Xbgfcpm__DUM_30 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_20 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_31 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_21 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_10 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_22 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_11 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__MB3_0 vdd vbn2 vdd vbp1 bgfcpm__MB3
Xbgfcpm__DUM_23 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_12 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__MB3_1 vdd vdd vbn2 vbp1 bgfcpm__MB3
Xbgfcpm__DUM_24 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_13 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__MB3_2 vdd vbn2 vdd vbp1 bgfcpm__MB3
Xbgfcpm__DUM_0 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_25 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_14 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__MB3_3 vdd vdd vbn2 vbp1 bgfcpm__MB3
Xbgfcpm__DUM_1 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_15 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_26 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_2 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_16 vdd vdd vdd vdd bgfcpm__DUM
Xbgfcpm__DUM_27 vdd vdd vdd vdd bgfcpm__DUM
.ends

.subckt bgfcnm__M4 a_100_n131# a_n100_n157# a_n158_n131# VSUBS
X0 a_100_n131# a_n100_n157# a_n158_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfcnm__M5 a_100_n131# a_n100_n157# a_n158_n131# VSUBS
X0 a_100_n131# a_n100_n157# a_n158_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfcnm__MB5 a_100_n131# a_n100_n157# a_n158_n131# VSUBS
X0 a_100_n131# a_n100_n157# a_n158_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfcnm__DUM a_100_n131# a_n100_n157# a_n158_n131# VSUBS
X0 a_100_n131# a_n100_n157# a_n158_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt bgfc__nmirr vbn1 out1n out1p vss
Xbgfcnm__M4_13 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M4_0 vss vbn1 out1n vss bgfcnm__M4
Xbgfcnm__M4_14 vss vbn1 out1n vss bgfcnm__M4
Xbgfcnm__M4_1 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M4_15 vss vbn1 out1n vss bgfcnm__M4
Xbgfcnm__M4_2 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M4_3 vss vbn1 out1n vss bgfcnm__M4
Xbgfcnm__M4_4 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M4_5 vss vbn1 out1n vss bgfcnm__M4
Xbgfcnm__M4_6 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M4_7 vss vbn1 out1n vss bgfcnm__M4
Xbgfcnm__M4_8 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M5_10 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__MB5_0 vbn1 vbn1 vss vss bgfcnm__MB5
Xbgfcnm__M4_9 vss vbn1 out1n vss bgfcnm__M4
Xbgfcnm__MB5_1 vss vbn1 vbn1 vss bgfcnm__MB5
Xbgfcnm__M5_11 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__M5_12 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__MB5_2 vss vbn1 vbn1 vss bgfcnm__MB5
Xbgfcnm__DUM_40 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_13 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__MB5_3 vbn1 vbn1 vss vss bgfcnm__MB5
Xbgfcnm__DUM_41 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_30 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_42 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_31 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_14 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__DUM_20 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_15 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__DUM_21 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_32 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_43 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_0 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_10 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_33 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_22 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_11 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_1 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_23 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_34 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_12 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_2 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_0 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__DUM_35 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_24 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_13 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_3 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_1 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__DUM_36 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_25 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_14 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_4 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_2 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__DUM_37 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_26 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_15 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_5 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_3 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__DUM_38 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_27 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_16 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_6 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_4 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__DUM_39 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_28 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_17 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_7 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_5 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__DUM_29 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_18 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_8 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_6 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__DUM_9 vss vss vss vss bgfcnm__DUM
Xbgfcnm__DUM_19 vss vss vss vss bgfcnm__DUM
Xbgfcnm__M5_7 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__M5_8 vss vbn1 out1p vss bgfcnm__M5
Xbgfcnm__M5_9 out1p vbn1 vss vss bgfcnm__M5
Xbgfcnm__M4_10 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M4_11 out1n vbn1 vss vss bgfcnm__M4
Xbgfcnm__M4_12 vss vbn1 out1n vss bgfcnm__M4
.ends

.subckt bgfccpt__DUM a_n458_n236# a_n400_n262# w_n494_n298# a_400_n236#
X0 a_400_n236# a_n400_n262# a_n458_n236# w_n494_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt bgfccpt__M11 a_n458_n236# a_n400_n262# w_n494_n298# a_400_n236#
X0 a_400_n236# a_n400_n262# a_n458_n236# w_n494_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt bgfccpt__M10 a_n458_n236# a_n400_n262# w_n494_n298# a_400_n236#
X0 a_400_n236# a_n400_n262# a_n458_n236# w_n494_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt bgfc__casp_top vdd nd11 nd10 mirr m1_458_30#
Xbgfccpt__DUM_7 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_8 mirr mirr m1_458_30# mirr bgfccpt__DUM
Xbgfccpt__M11_0 vdd mirr m1_458_30# nd11 bgfccpt__M11
Xbgfccpt__DUM_9 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__M11_1 nd11 mirr m1_458_30# vdd bgfccpt__M11
Xbgfccpt__DUM_20 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__M11_2 vdd mirr m1_458_30# nd11 bgfccpt__M11
Xbgfccpt__DUM_21 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_10 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__M11_3 nd11 mirr m1_458_30# vdd bgfccpt__M11
Xbgfccpt__DUM_22 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_11 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__M11_4 nd11 mirr m1_458_30# vdd bgfccpt__M11
Xbgfccpt__DUM_12 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_23 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__M11_5 vdd mirr m1_458_30# nd11 bgfccpt__M11
Xbgfccpt__DUM_13 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__M11_6 vdd mirr m1_458_30# nd11 bgfccpt__M11
Xbgfccpt__DUM_14 mirr mirr m1_458_30# mirr bgfccpt__DUM
Xbgfccpt__M11_7 nd11 mirr m1_458_30# vdd bgfccpt__M11
Xbgfccpt__DUM_15 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_16 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_17 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_18 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_19 mirr mirr m1_458_30# mirr bgfccpt__DUM
Xbgfccpt__M10_0 vdd mirr m1_458_30# nd10 bgfccpt__M10
Xbgfccpt__M10_1 nd10 mirr m1_458_30# vdd bgfccpt__M10
Xbgfccpt__M10_2 nd10 mirr m1_458_30# vdd bgfccpt__M10
Xbgfccpt__M10_3 nd10 mirr m1_458_30# vdd bgfccpt__M10
Xbgfccpt__M10_4 vdd mirr m1_458_30# nd10 bgfccpt__M10
Xbgfccpt__M10_5 nd10 mirr m1_458_30# vdd bgfccpt__M10
Xbgfccpt__M10_6 vdd mirr m1_458_30# nd10 bgfccpt__M10
Xbgfccpt__M10_7 vdd mirr m1_458_30# nd10 bgfccpt__M10
Xbgfccpt__DUM_0 mirr mirr m1_458_30# mirr bgfccpt__DUM
Xbgfccpt__DUM_1 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_2 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_3 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_4 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_5 vdd vdd m1_458_30# vdd bgfccpt__DUM
Xbgfccpt__DUM_6 vdd vdd m1_458_30# vdd bgfccpt__DUM
.ends

.subckt bgfccnt__M6 a_400_n131# a_n400_n157# a_n458_n131# VSUBS
X0 a_400_n131# a_n400_n157# a_n458_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
.ends

.subckt bgfccnt__DUM a_400_n131# a_n400_n157# a_n458_n131# VSUBS
X0 a_400_n131# a_n400_n157# a_n458_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
.ends

.subckt bgfccnt__M7 a_400_n131# a_n400_n157# a_n458_n131# VSUBS
X0 a_400_n131# a_n400_n157# a_n458_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
.ends

.subckt bgfccnt__MB4 a_400_n131# a_n400_n157# a_n458_n131# VSUBS
X0 a_400_n131# a_n400_n157# a_n458_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=4
.ends

.subckt bgfc__casn_top vbn2 vbn1 mirr out1n out1p out VSUBS
Xbgfccnt__M6_0 mirr vbn2 out1n VSUBS bgfccnt__M6
Xbgfccnt__M6_1 out1n vbn2 mirr VSUBS bgfccnt__M6
Xbgfccnt__M6_2 out1n vbn2 mirr VSUBS bgfccnt__M6
Xbgfccnt__M6_3 mirr vbn2 out1n VSUBS bgfccnt__M6
Xbgfccnt__M6_4 out1n vbn2 mirr VSUBS bgfccnt__M6
Xbgfccnt__DUM_0 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__M6_5 mirr vbn2 out1n VSUBS bgfccnt__M6
Xbgfccnt__DUM_1 vbn2 vbn2 vbn2 VSUBS bgfccnt__DUM
Xbgfccnt__M6_6 out1n vbn2 mirr VSUBS bgfccnt__M6
Xbgfccnt__DUM_2 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__M6_7 mirr vbn2 out1n VSUBS bgfccnt__M6
Xbgfccnt__DUM_3 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_4 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_5 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_6 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_7 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_8 vbn2 vbn2 vbn2 VSUBS bgfccnt__DUM
Xbgfccnt__DUM_9 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__M7_0 out vbn2 out1p VSUBS bgfccnt__M7
Xbgfccnt__M7_1 out1p vbn2 out VSUBS bgfccnt__M7
Xbgfccnt__M7_2 out1p vbn2 out VSUBS bgfccnt__M7
Xbgfccnt__DUM_20 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__MB4_0 vbn1 vbn2 vbn2 VSUBS bgfccnt__MB4
Xbgfccnt__M7_3 out vbn2 out1p VSUBS bgfccnt__M7
Xbgfccnt__DUM_10 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_21 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__MB4_1 vbn1 vbn2 vbn2 VSUBS bgfccnt__MB4
Xbgfccnt__M7_4 out vbn2 out1p VSUBS bgfccnt__M7
Xbgfccnt__DUM_11 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_22 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__MB4_2 vbn2 vbn2 vbn1 VSUBS bgfccnt__MB4
Xbgfccnt__M7_5 out1p vbn2 out VSUBS bgfccnt__M7
Xbgfccnt__DUM_12 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_23 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__MB4_3 vbn2 vbn2 vbn1 VSUBS bgfccnt__MB4
Xbgfccnt__M7_6 out1p vbn2 out VSUBS bgfccnt__M7
Xbgfccnt__DUM_13 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_24 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__M7_7 out vbn2 out1p VSUBS bgfccnt__M7
Xbgfccnt__DUM_14 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_25 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_26 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_15 vbn2 vbn2 vbn2 VSUBS bgfccnt__DUM
Xbgfccnt__DUM_16 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_27 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_17 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_18 VSUBS VSUBS VSUBS VSUBS bgfccnt__DUM
Xbgfccnt__DUM_19 vbn2 vbn2 vbn2 VSUBS bgfccnt__DUM
.ends

.subckt bgfcdpp__M3 w_n194_n498# a_100_n436# a_n158_n436# a_n100_n462#
X0 a_100_n436# a_n100_n462# a_n158_n436# w_n194_n498# sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt bgfcdpp__M2 w_n194_n498# a_100_n436# a_n158_n436# a_n100_n462#
X0 a_100_n436# a_n100_n462# a_n158_n436# w_n194_n498# sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt bgfcdpp__DUM w_n194_n498# a_100_n436# a_n158_n436# a_n100_n462#
X0 a_100_n436# a_n100_n462# a_n158_n436# w_n194_n498# sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt bgfc__diffpair_p inp inn diff out1p out1n vdd
Xbgfcdpp__M3_0 vdd diff out1p inn bgfcdpp__M3
Xbgfcdpp__M3_1 vdd out1p diff inn bgfcdpp__M3
Xbgfcdpp__M3_2 vdd diff out1p inn bgfcdpp__M3
Xbgfcdpp__M3_3 vdd out1p diff inn bgfcdpp__M3
Xbgfcdpp__M3_4 vdd diff out1p inn bgfcdpp__M3
Xbgfcdpp__M3_5 vdd out1p diff inn bgfcdpp__M3
Xbgfcdpp__M3_6 vdd diff out1p inn bgfcdpp__M3
Xbgfcdpp__M3_7 vdd out1p diff inn bgfcdpp__M3
Xbgfcdpp__M2_0 vdd diff out1n inp bgfcdpp__M2
Xbgfcdpp__M2_1 vdd out1n diff inp bgfcdpp__M2
Xbgfcdpp__M2_2 vdd diff out1n inp bgfcdpp__M2
Xbgfcdpp__M2_3 vdd out1n diff inp bgfcdpp__M2
Xbgfcdpp__M2_4 vdd diff out1n inp bgfcdpp__M2
Xbgfcdpp__M2_5 vdd out1n diff inp bgfcdpp__M2
Xbgfcdpp__M2_6 vdd out1n diff inp bgfcdpp__M2
Xbgfcdpp__M2_7 vdd diff out1n inp bgfcdpp__M2
Xbgfcdpp__DUM_0 vdd diff diff diff bgfcdpp__DUM
Xbgfcdpp__DUM_1 vdd diff diff diff bgfcdpp__DUM
Xbgfcdpp__DUM_2 vdd diff diff diff bgfcdpp__DUM
Xbgfcdpp__DUM_3 vdd diff diff diff bgfcdpp__DUM
.ends

.subckt bgfccpb__M8 a_n458_n236# a_n400_n262# w_n494_n298# a_400_n236#
X0 a_400_n236# a_n400_n262# a_n458_n236# w_n494_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt bgfccpb__M9 a_n458_n236# a_n400_n262# w_n494_n298# a_400_n236#
X0 a_400_n236# a_n400_n262# a_n458_n236# w_n494_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt bgfccpb__DUM a_n458_n236# a_n400_n262# w_n494_n298# a_400_n236#
X0 a_400_n236# a_n400_n262# a_n458_n236# w_n494_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt bgfccpb__MB1 a_n458_n236# a_n400_n262# w_n494_n298# a_400_n236#
X0 a_400_n236# a_n400_n262# a_n458_n236# w_n494_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
.ends

.subckt bgfc__casp_bot nd11 nd10 mirr bias vbp1 out m1_458_17#
Xbgfccpb__M8_0 mirr bias m1_458_17# nd10 bgfccpb__M8
Xbgfccpb__M8_1 nd10 bias m1_458_17# mirr bgfccpb__M8
Xbgfccpb__M8_2 mirr bias m1_458_17# nd10 bgfccpb__M8
Xbgfccpb__M8_3 nd10 bias m1_458_17# mirr bgfccpb__M8
Xbgfccpb__M8_4 nd10 bias m1_458_17# mirr bgfccpb__M8
Xbgfccpb__M8_5 mirr bias m1_458_17# nd10 bgfccpb__M8
Xbgfccpb__M8_6 nd10 bias m1_458_17# mirr bgfccpb__M8
Xbgfccpb__M8_7 mirr bias m1_458_17# nd10 bgfccpb__M8
Xbgfccpb__M9_0 out bias m1_458_17# nd11 bgfccpb__M9
Xbgfccpb__M9_1 nd11 bias m1_458_17# out bgfccpb__M9
Xbgfccpb__DUM_0 bias bias m1_458_17# bias bgfccpb__DUM
Xbgfccpb__M9_2 nd11 bias m1_458_17# out bgfccpb__M9
Xbgfccpb__MB1_0 vbp1 bias m1_458_17# bias bgfccpb__MB1
Xbgfccpb__M9_3 out bias m1_458_17# nd11 bgfccpb__M9
Xbgfccpb__DUM_1 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__MB1_1 vbp1 bias m1_458_17# bias bgfccpb__MB1
Xbgfccpb__DUM_2 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__M9_4 nd11 bias m1_458_17# out bgfccpb__M9
Xbgfccpb__MB1_2 bias bias m1_458_17# vbp1 bgfccpb__MB1
Xbgfccpb__M9_5 out bias m1_458_17# nd11 bgfccpb__M9
Xbgfccpb__DUM_3 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_20 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__MB1_3 bias bias m1_458_17# vbp1 bgfccpb__MB1
Xbgfccpb__DUM_4 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__M9_6 nd11 bias m1_458_17# out bgfccpb__M9
Xbgfccpb__DUM_21 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_10 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__M9_7 out bias m1_458_17# nd11 bgfccpb__M9
Xbgfccpb__DUM_5 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_22 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_11 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_6 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_23 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_12 bias bias m1_458_17# bias bgfccpb__DUM
Xbgfccpb__DUM_7 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_24 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_13 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_8 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_14 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_25 bias bias m1_458_17# bias bgfccpb__DUM
Xbgfccpb__DUM_9 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_26 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_15 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_16 bias bias m1_458_17# bias bgfccpb__DUM
Xbgfccpb__DUM_27 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_17 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_18 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
Xbgfccpb__DUM_19 m1_458_17# m1_458_17# m1_458_17# m1_458_17# bgfccpb__DUM
.ends

.subckt bg__se_folded_cascode_p vbn1 vbp1 diff out1p out1n mirr vbn2 nd10 nd11 out
+ vdd bias vsub inp inn vss
Xbgfc__pmirr_0 vbp1 diff vbn2 vdd bgfc__pmirr
Xbgfc__nmirr_0 vbn1 out1n out1p vss bgfc__nmirr
Xbgfc__casp_top_0 vdd nd11 nd10 mirr vdd bgfc__casp_top
Xbgfc__casn_top_0 vbn2 vbn1 mirr out1n out1p out vss bgfc__casn_top
Xbgfc__diffpair_p_0 inp inn diff out1p out1n vdd bgfc__diffpair_p
Xbgfc__casp_bot_0 nd11 nd10 mirr bias vbp1 out vdd bgfc__casp_bot
.ends

.subckt bandgap_cw vbg trim[15] trim[13] trim[11] trim[9] trim[7] trim[5] trim[3]
+ trim[1] trim[0] trim[2] trim[4] trim[6] trim[8] trim[10] trim[12] trim[14] bias
+ vdd vsub vss
Xbg__cap_3 bg__se_folded_cascode_p_0/out vss bg__cap
Xbg__cap_4 bg__se_folded_cascode_p_0/out vss bg__cap
Xbg__res_0 m1_32787_8825# m1_32015_12378# m1_35489_12378# m1_30085_12378# m1_33559_12378#
+ m1_30857_8825# m1_35103_12378# m1_31243_9043# m1_30085_12378# m1_29699_9043# m1_29699_9043#
+ m2_32390_12378# m1_35103_12378# m1_28541_12378# m1_34717_9043# m1_30471_12378# m1_31629_12378#
+ m1_34717_9043# m1_33977_7455# m1_28927_12378# bg__se_folded_cascode_p_0/inp m1_32787_8825#
+ m1_33173_9043# m1_33559_12378# m1_34331_8825# m1_33945_12378# m1_29313_8825# bg__se_folded_cascode_p_0/inp
+ m1_31629_12378# m1_35489_12378# bg__pnp_group_0/eu m1_30471_12378# m1_32015_12378#
+ m1_33945_12378# m1_34331_8825# m1_28927_12378# m1_31243_9043# vbg m1_30857_8825#
+ m1_28541_12378# m1_29313_8825# vss m1_33173_9043# bg__res
Xbg__cap_5 bg__se_folded_cascode_p_0/out vss bg__cap
Xbg__cap_6 bg__se_folded_cascode_p_0/out vss bg__cap
Xbg__cap_7 bg__se_folded_cascode_p_0/out vss bg__cap
Xbg__cap_8 m4_36893_6523# vss bg__cap
Xbg__trim_0 trim[7] trim[10] trim[8] trim[1] bg__pnp_group_0/eg trim[14] trim[6] trim[5]
+ trim[4] bg__pnp_group_0/eg bg__pnp_group_0/eg trim[11] trim[15] trim[2] m2_32390_12378#
+ trim[9] trim[3] trim[12] trim[0] vss trim[13] bg__trim
Xbg__cap_9 m4_36893_6523# vss bg__cap
Xbg__startup_0 vbg vss vss vdd vdd vdd m4_36893_6523# m4_36893_6523# bg__se_folded_cascode_p_0/out
+ vss bg__startup
Xbg__M1_M2_0 vbg bg__se_folded_cascode_p_0/out vdd m1_33977_7455# bg__se_folded_cascode_p_0/out
+ vdd vdd bg__se_folded_cascode_p_0/out vdd bg__se_folded_cascode_p_0/out bg__M1_M2
Xbg__pnp_group_0 bg__pnp_group_0/eg bg__pnp_group_0/eu vdd vss bg__pnp_group
Xbg__cap_10 m4_36893_6523# vss bg__cap
Xbg__se_folded_cascode_p_0 bg__se_folded_cascode_p_0/vbn1 bg__se_folded_cascode_p_0/vbp1
+ bg__se_folded_cascode_p_0/diff bg__se_folded_cascode_p_0/out1p bg__se_folded_cascode_p_0/out1n
+ bg__se_folded_cascode_p_0/mirr bg__se_folded_cascode_p_0/vbn2 bg__se_folded_cascode_p_0/nd10
+ bg__se_folded_cascode_p_0/nd11 bg__se_folded_cascode_p_0/out vdd bias vsub bg__se_folded_cascode_p_0/inp
+ bg__pnp_group_0/eu vss bg__se_folded_cascode_p
Xbg__cap_0 bg__se_folded_cascode_p_0/out vss bg__cap
Xbg__cap_1 bg__se_folded_cascode_p_0/out vss bg__cap
Xbg__cap_2 bg__se_folded_cascode_p_0/out vss bg__cap
.ends

.subckt sky130_cw_ip__bandgap_nobias trim[0] trim[4] trim[6] trim[10] trim[12] trim[14]
+ trim[15] trim[13] trim[11] trim[7] trim[5] trim[3] trim[1] trim[2] vsub bias vbg
+ trim[9] trim[8] vdd vss
Xbandgap_cw_0 vbg trim[15] trim[13] trim[11] trim[9] trim[7] trim[5] trim[3] trim[1]
+ trim[0] trim[2] trim[4] trim[6] trim[8] trim[10] trim[12] trim[14] bias vdd vsub
+ vss bandgap_cw
.ends

.subckt frigate_analog gpio5_4 gpio5_5 gpio5_6 gpio5_7 gpio6_0 gpio6_1 gpio6_2 gpio6_3
+ left_vref gpio6_4 gpio6_5 gpio6_6 gpio6_7 adc_refl_to_gpio6_7[1] adc_refl_to_gpio6_7[0]
+ adc_refh_to_gpio6_6[1] adc_refh_to_gpio6_6[0] adc1_to_gpio6_5[1] adc1_to_gpio6_5[0]
+ adc0_to_gpio6_4[1] adc0_to_gpio6_4[0] comp_p_to_gpio6_2[1] comp_p_to_gpio6_2[0]
+ comp_n_to_gpio6_3[1] comp_n_to_gpio6_3[0] ulpcomp_n_to_gpio6_1[1] ulpcomp_n_to_gpio6_1[0]
+ ulpcomp_p_to_gpio6_0[1] ulpcomp_p_to_gpio6_0[0] left_instramp_n_to_gpio5_7[1] left_instramp_n_to_gpio5_7[0]
+ left_instramp_p_to_gpio5_6[1] left_instramp_p_to_gpio5_6[0] left_lp_opamp_n_to_gpio5_5[1]
+ left_lp_opamp_n_to_gpio5_5[0] left_lp_opamp_p_to_gpio5_4[1] left_lp_opamp_p_to_gpio5_4[0]
+ left_hgbw_opamp_n_to_gpio5_3[1] left_hgbw_opamp_n_to_gpio5_3[0] left_hgbw_opamp_p_to_gpio5_2[1]
+ left_hgbw_opamp_p_to_gpio5_2[0] right_hgbw_opamp_n_to_gpio5_1[1] right_hgbw_opamp_n_to_gpio5_1[0]
+ right_hgbw_opamp_p_to_gpio5_0[1] right_hgbw_opamp_p_to_gpio5_0[0] right_lp_opamp_to_gpio4_7[1]
+ right_lp_opamp_to_gpio4_7[0] right_hgbw_opamp_to_gpio4_6[1] right_hgbw_opamp_to_gpio4_6[0]
+ left_hgbw_opamp_to_gpio4_5[1] left_hgbw_opamp_to_gpio4_5[0] left_instramp_to_gpio4_4[1]
+ left_instramp_to_gpio4_4[0] right_lp_opamp_to_gpio4_3[1] right_lp_opamp_to_gpio4_3[0]
+ right_hgbw_opamp_to_gpio4_2[1] right_hgbw_opamp_to_gpio4_2[0] left_hgbw_opamp_to_gpio4_1[1]
+ left_hgbw_opamp_to_gpio4_1[0] left_lp_opamp_to_gpio4_0[1] left_lp_opamp_to_gpio4_0[0]
+ left_instramp_to_ulpcomp_p[1] left_instramp_to_ulpcomp_p[0] left_instramp_to_comp_p[1]
+ left_instramp_to_comp_p[0] left_instramp_to_adc0[1] left_instramp_to_adc0[0] left_instramp_to_analog1[1]
+ left_instramp_to_analog1[0] left_instramp_to_amuxbusB[1] left_instramp_to_amuxbusB[0]
+ left_instramp_n_to_analog1 left_instramp_n_to_amuxbusB right_lp_opamp_to_ulpcomp_p[1]
+ right_lp_opamp_to_ulpcomp_p[0] right_lp_opamp_to_comp_p[1] right_lp_opamp_to_comp_p[0]
+ right_lp_opamp_to_adc0[1] right_lp_opamp_to_adc0[0] right_hgbw_opamp_to_ulpcomp_n[1]
+ right_hgbw_opamp_to_ulpcomp_n[0] right_hgbw_opamp_to_comp_n[1] right_hgbw_opamp_to_comp_n[0]
+ right_hgbw_opamp_to_adc1[1] right_hgbw_opamp_to_adc1[0] right_instramp_to_ulpcomp_n[1]
+ right_instramp_to_ulpcomp_n[0] right_instramp_to_comp_n[1] right_instramp_to_comp_n[0]
+ right_instramp_to_adc1[1] right_instramp_to_adc1[0] left_instramp_p_to_analog0 left_instramp_p_to_amuxbusA
+ left_hgbw_opamp_to_ulpcomp_p[1] left_hgbw_opamp_to_ulpcomp_p[0] left_hgbw_opamp_to_comp_p[1]
+ left_hgbw_opamp_to_comp_p[0] left_hgbw_opamp_to_adc0[1] left_hgbw_opamp_to_adc0[0]
+ left_hgbw_opamp_to_analog1[1] left_hgbw_opamp_to_analog1[0] left_hgbw_opamp_to_amuxbusB[1]
+ left_hgbw_opamp_to_amuxbusB[0] left_hgbw_opamp_p_to_dac0 left_hgbw_opamp_p_to_analog0
+ left_hgbw_opamp_p_to_amuxbusA left_instramp_p_to_left_rheostat1_out left_hgbw_opamp_n_to_dac1
+ left_hgbw_opamp_n_to_analog1 left_hgbw_opamp_n_to_amuxbusB left_instramp_n_to_left_rheostat1_out
+ left_hgbw_opamp_n_to_rheostat_tap left_lp_opamp_to_ulpcomp_n[1] left_lp_opamp_to_ulpcomp_n[0]
+ left_lp_opamp_to_comp_n[1] left_lp_opamp_to_comp_n[0] left_lp_opamp_to_adc1[1] left_lp_opamp_to_adc1[0]
+ left_lp_opamp_to_analog0[1] left_lp_opamp_to_analog0[0] left_lp_opamp_to_amuxbusA[1]
+ left_lp_opamp_to_amuxbusA[0] left_lp_opamp_p_to_dac0 left_lp_opamp_p_to_analog0
+ left_lp_opamp_p_to_amuxbusA right_instramp_p_to_left_rheostat2_out left_lp_opamp_n_to_dac1
+ left_lp_opamp_n_to_analog1 left_lp_opamp_n_to_amuxbusB right_instramp_n_to_left_rheostat2_out
+ left_lp_opamp_n_to_rheostat_tap adc0_to_dac0 adc0_to_analog1 adc1_to_dac1 adc1_to_analog0
+ vdda1_pwr_good vccd1_pwr_good vdda2_pwr_good vccd2_pwr_good audiodac_in adc0_dac_val[15]
+ adc0_comp_out adc0_hold adc0_reset adc1_dac_val[15] adc1_comp_out adc1_hold adc1_reset
+ tempsense_ena rdac0_ena rdac0_value[11] rdac0_value[10] rdac0_value[9] rdac0_value[8]
+ rdac0_value[7] rdac0_value[6] rdac0_value[5] rdac0_value[4] rdac0_value[3] rdac0_value[2]
+ rdac0_value[1] rdac0_value[0] rdac1_ena rdac1_value[11] rdac1_value[10] rdac1_value[9]
+ rdac1_value[8] rdac1_value[7] rdac1_value[6] rdac1_value[5] rdac1_value[4] rdac1_value[3]
+ rdac1_value[2] rdac1_value[1] rdac1_value[0] adc0_ena adc1_ena left_instramp_ena
+ left_instramp_G1[4] left_instramp_G1[3] left_instramp_G1[2] left_instramp_G1[1]
+ left_instramp_G1[0] left_instramp_G2[4] left_instramp_G2[3] left_instramp_G2[2]
+ left_instramp_G2[1] left_instramp_G2[0] left_hgbw_opamp_ena left_lp_opamp_ena left_rheostat1_b[7]
+ left_rheostat1_b[6] left_rheostat1_b[5] left_rheostat1_b[4] left_rheostat1_b[3]
+ left_rheostat1_b[2] left_rheostat1_b[1] left_rheostat1_b[0] left_rheostat2_b[7]
+ left_rheostat2_b[6] left_rheostat2_b[5] left_rheostat2_b[4] left_rheostat2_b[3]
+ left_rheostat2_b[2] left_rheostat2_b[1] left_rheostat2_b[0] analog0_connect[1] analog0_connect[0]
+ analog1_connect[1] analog1_connect[0] user_voutref user_vinref user_left_vref user_right_vref
+ user_tempsense user_dac0 user_dac1 user_vbgtc user_vbgsc user_adc0 user_adc1 user_comp_n
+ user_comp_p user_ulpcomp_n user_ulpcomp_p user_gpio4_7_analog user_gpio4_6_analog
+ user_gpio4_5_analog user_gpio4_4_analog user_gpio4_3_analog user_gpio4_2_analog
+ user_gpio4_1_analog user_gpio4_0_analog user_gpio3_7_analog user_gpio3_6_analog
+ user_gpio3_5_analog user_gpio3_4_analog user_gpio3_3_analog user_gpio3_2_analog
+ user_gpio3_1_analog user_gpio3_0_analog comp_out ulpcomp_out overvoltage_out comp_ena
+ comp_trim[5] comp_trim[4] comp_trim[3] comp_trim[2] comp_trim[1] comp_trim[0] comp_hyst[1]
+ comp_hyst[0] ulpcomp_ena ulpcomp_clk bandgap_ena bandgap_trim[15] bandgap_trim[14]
+ bandgap_trim[13] bandgap_trim[12] bandgap_trim[11] bandgap_trim[10] bandgap_trim[9]
+ bandgap_trim[8] bandgap_trim[7] bandgap_trim[6] bandgap_trim[5] bandgap_trim[4]
+ bandgap_trim[3] bandgap_trim[2] bandgap_trim[1] bandgap_trim[0] ldo_ena ibias_ena
+ ibias_src_ena[23] ibias_src_ena[22] ibias_src_ena[21] ibias_src_ena[20] ibias_src_ena[19]
+ ibias_src_ena[18] ibias_src_ena[17] ibias_src_ena[16] ibias_src_ena[15] ibias_src_ena[14]
+ ibias_src_ena[13] ibias_src_ena[12] ibias_src_ena[11] ibias_src_ena[10] ibias_src_ena[9]
+ ibias_src_ena[8] ibias_src_ena[7] ibias_src_ena[6] ibias_src_ena[5] ibias_src_ena[4]
+ ibias_src_ena[3] ibias_src_ena[2] ibias_src_ena[1] ibias_src_ena[0] ibias_snk_ena[3]
+ ibias_snk_ena[2] ibias_snk_ena[1] ibias_snk_ena[0] ibias_ref_select overvoltage_ena
+ overvoltage_trim[3] overvoltage_trim[2] overvoltage_trim[1] overvoltage_trim[0]
+ idac_value[11] idac_value[10] idac_value[9] idac_value[8] idac_value[7] idac_value[6]
+ idac_value[5] idac_value[4] idac_value[3] idac_value[2] idac_value[1] idac_value[0]
+ idac_ena right_instramp_ena right_instramp_G1[4] right_instramp_G1[3] right_instramp_G1[2]
+ right_instramp_G1[1] right_instramp_G1[0] right_instramp_G2[4] right_instramp_G2[3]
+ right_instramp_G2[2] right_instramp_G2[1] right_instramp_G2[0] right_hgbw_opamp_ena
+ right_lp_opamp_ena right_rheostat1_b[7] right_rheostat1_b[6] right_rheostat1_b[5]
+ right_rheostat1_b[4] right_rheostat1_b[3] right_rheostat1_b[2] right_rheostat1_b[1]
+ right_rheostat1_b[0] right_rheostat2_b[7] right_rheostat2_b[6] right_rheostat2_b[5]
+ right_rheostat2_b[4] right_rheostat2_b[3] right_rheostat2_b[2] right_rheostat2_b[1]
+ right_rheostat2_b[0] por porb porb_h[1] user_to_comp_n[1] user_to_comp_n[0] user_to_comp_p[1]
+ user_to_comp_p[0] user_to_ulpcomp_n[1] user_to_ulpcomp_n[0] user_to_ulpcomp_p[1]
+ user_to_ulpcomp_p[0] user_to_adc0[1] user_to_adc0[0] user_to_adc1[1] user_to_adc1[0]
+ dac0_to_user dac1_to_user tempsense_to_user right_vref_to_user left_vref_to_user
+ vinref_to_user voutref_to_user vbgtc_to_user vbgsc_to_user sio0_connect[1] sio0_connect[0]
+ sio1_connect[1] sio1_connect[0] comp_p_to_dac0 comp_p_to_analog1 comp_p_to_sio0
+ comp_p_to_vbgtc comp_p_to_tempsense comp_p_to_left_vref comp_p_to_voutref comp_n_to_dac1
+ comp_n_to_analog0 comp_n_to_sio1 comp_n_to_vbgsc comp_n_to_right_vref comp_n_to_vinref
+ ulpcomp_p_to_dac0 ulpcomp_p_to_analog1 ulpcomp_p_to_sio0 ulpcomp_p_to_vbgtc ulpcomp_p_to_tempsense
+ ulpcomp_p_to_left_vref ulpcomp_p_to_voutref ulpcomp_n_to_dac1 ulpcomp_n_to_analog0
+ ulpcomp_n_to_sio1 ulpcomp_n_to_vbgsc ulpcomp_n_to_right_vref ulpcomp_n_to_vinref
+ left_instramp_n_to_sio1 left_instramp_n_to_right_vref left_instramp_n_to_vinref
+ left_instramp_p_to_sio0 left_instramp_p_to_tempsense left_instramp_p_to_left_vref
+ left_instramp_p_to_voutref left_hgbw_opamp_p_to_sio0 left_hgbw_opamp_p_to_tempsense
+ left_hgbw_opamp_p_to_left_vref left_hgbw_opamp_p_to_voutref left_lp_opamp_p_to_sio0
+ left_lp_opamp_p_to_left_vref left_lp_opamp_p_to_voutref left_hgbw_opamp_n_to_sio1
+ left_hgbw_opamp_n_to_vbgtc left_hgbw_opamp_n_to_right_vref left_hgbw_opamp_n_to_vinref
+ left_lp_opamp_n_to_sio1 left_lp_opamp_n_to_vbgsc left_lp_opamp_n_to_right_vref left_lp_opamp_n_to_vinref
+ adc0_to_vbgtc adc0_to_tempsense adc0_to_left_vref adc0_to_voutref adc1_to_vbgsc
+ adc1_to_right_vref adc1_to_vinref right_lp_opamp_to_analog1[1] right_lp_opamp_to_analog1[0]
+ right_lp_opamp_to_amuxbusB[1] right_lp_opamp_to_amuxbusB[0] right_lp_opamp_p_to_dac0
+ right_lp_opamp_p_to_analog0 right_lp_opamp_p_to_amuxbusA left_instramp_p_to_right_rheostat2_out
+ right_lp_opamp_p_to_sio0 right_lp_opamp_p_to_tempsense right_lp_opamp_p_to_left_vref
+ right_lp_opamp_p_to_voutref right_lp_opamp_n_to_dac1 right_lp_opamp_n_to_analog1
+ right_lp_opamp_n_to_amuxbusB left_instramp_n_to_right_rheostat2_out right_lp_opamp_n_to_rheostat_tap
+ right_lp_opamp_n_to_sio1 right_lp_opamp_n_to_vbgtc right_lp_opamp_n_to_right_vref
+ right_lp_opamp_n_to_vinref right_hgbw_opamp_to_analog0[1] right_hgbw_opamp_to_analog0[0]
+ right_hgbw_opamp_to_amuxbusA[1] right_hgbw_opamp_to_amuxbusA[0] right_hgbw_opamp_p_to_dac0
+ right_hgbw_opamp_p_to_analog0 right_hgbw_opamp_p_to_amuxbusA right_instramp_p_to_right_rheostat1_out
+ right_hgbw_opamp_p_to_sio0 right_hgbw_opamp_p_to_left_vref right_hgbw_opamp_p_to_voutref
+ right_hgbw_opamp_n_to_dac1 right_hgbw_opamp_n_to_analog1 right_hgbw_opamp_n_to_amuxbusB
+ right_instramp_n_to_right_rheostat1_out right_hgbw_opamp_n_to_rheostat_tap right_hgbw_opamp_n_to_sio1
+ right_hgbw_opamp_n_to_vbgsc right_hgbw_opamp_n_to_right_vref right_hgbw_opamp_n_to_vinref
+ right_instramp_to_analog0[1] right_instramp_to_analog0[0] right_instramp_to_amuxbusA[1]
+ right_instramp_to_amuxbusA[0] right_instramp_n_to_analog1 right_instramp_n_to_amuxbusB
+ right_instramp_n_to_sio1 right_instramp_n_to_right_vref right_instramp_n_to_vinref
+ right_instramp_p_to_analog0 right_instramp_p_to_amuxbusA right_instramp_p_to_tempsense
+ right_instramp_p_to_left_vref right_instramp_p_to_voutref right_lp_opamp_to_gpio3_7[1]
+ right_lp_opamp_to_gpio3_7[0] right_hgbw_opamp_to_gpio3_6[1] right_hgbw_opamp_to_gpio3_6[0]
+ left_hgbw_opamp_to_gpio3_5[1] left_hgbw_opamp_to_gpio3_5[0] left_lp_opamp_to_gpio3_4[1]
+ left_lp_opamp_to_gpio3_4[0] right_lp_opamp_to_gpio3_3[1] right_lp_opamp_to_gpio3_3[0]
+ right_hgbw_opamp_to_gpio3_2[1] right_hgbw_opamp_to_gpio3_2[0] left_hgbw_opamp_to_gpio3_1[1]
+ left_hgbw_opamp_to_gpio3_1[0] right_instramp_to_gpio3_0[1] right_instramp_to_gpio3_0[0]
+ right_instramp_p_to_gpio2_7[1] right_instramp_p_to_gpio2_7[0] right_instramp_n_to_gpio2_6[1]
+ right_instramp_n_to_gpio2_6[0] right_lp_opamp_p_to_gpio2_5[1] right_lp_opamp_p_to_gpio2_5[0]
+ right_lp_opamp_n_to_gpio2_4[1] right_lp_opamp_n_to_gpio2_4[0] right_hgbw_opamp_p_to_gpio2_3[1]
+ right_hgbw_opamp_p_to_gpio2_3[0] right_hgbw_opamp_n_to_gpio2_2[1] right_hgbw_opamp_n_to_gpio2_2[0]
+ left_hgbw_opamp_p_to_gpio2_1[1] left_hgbw_opamp_p_to_gpio2_1[0] left_hgbw_opamp_n_to_gpio2_0[1]
+ left_hgbw_opamp_n_to_gpio2_0[0] ulpcomp_p_to_gpio1_7[1] ulpcomp_p_to_gpio1_7[0]
+ ulpcomp_n_to_gpio1_6[1] ulpcomp_n_to_gpio1_6[0] comp_p_to_gpio1_5[1] comp_p_to_gpio1_5[0]
+ comp_n_to_gpio1_4[1] comp_n_to_gpio1_4[0] adc0_to_gpio1_3[1] adc0_to_gpio1_3[0]
+ idac_to_gpio1_3[1] idac_to_gpio1_3[0] ibias_test_to_gpio1_2[1] ibias_test_to_gpio1_2[0]
+ idac_to_gpio1_2[1] idac_to_gpio1_2[0] adc1_to_gpio1_2[1] adc1_to_gpio1_2[0] dac_refh_to_gpio1_1[1]
+ dac_refh_to_gpio1_1[0] vbg_test_to_gpio1_1[1] vbg_test_to_gpio1_1[0] dac_refl_to_gpio1_0[1]
+ dac_refl_to_gpio1_0[0] ibias_lsxo ibias_hsxo sio0 sio1 voutref vinref vbg gpio2_3
+ gpio2_2 gpio2_1 gpio2_0 gpio1_7 gpio1_6 gpio1_5 gpio1_4 right_vref gpio1_3 gpio1_2
+ gpio1_1 gpio1_0 gpio5_3 gpio5_2 gpio5_1 gpio5_0 gpio4_7 gpio4_6 gpio4_5 gpio4_4
+ gpio4_3 gpio4_2 gpio4_1 gpio4_0 analog1 analog0 amuxbus_b_n amuxbus_a_n gpio3_7
+ gpio3_6 gpio3_5 gpio3_4 gpio3_3 gpio3_2 gpio3_1 gpio3_0 gpio2_4 gpio2_5 gpio2_6
+ gpio2_7 vdda2 vssa2 vccd2 vssd2 vssd1 vccd1 vssa1 vdda1 user_ibias50 user_ibias100
+ vdda0 vssa0 audiodac_inb audiodac_outb_to_analog0[1] audiodac_out_to_analog1[1]
+ bandgap_sel ldo_ref_sel tempsense_sel vddio vssio vssd0 vccd0 right_instramp_p_to_sio0
+ brownout_ena brownout_vtrip[2] brownout_vtrip[1] brownout_vtrip[0] brownout_otrip[2]
+ brownout_otrip[1] brownout_otrip[0] brownout_isrc_sel brownout_oneshot brownout_rc_ena
+ brownout_rc_dis brownout_vunder brownout_timeout brownout_filt brownout_unfilt dac1_to_analog0
+ dac0_to_analog1 adc1_dac_val[14] adc1_dac_val[13] adc1_dac_val[12] adc1_dac_val[11]
+ adc1_dac_val[10] adc1_dac_val[9] adc1_dac_val[8] adc1_dac_val[7] adc1_dac_val[6]
+ adc1_dac_val[5] adc1_dac_val[4] adc1_dac_val[3] adc1_dac_val[2] adc1_dac_val[1]
+ adc1_dac_val[0] adc0_dac_val[14] adc0_dac_val[13] adc0_dac_val[12] adc0_dac_val[11]
+ adc0_dac_val[10] adc0_dac_val[9] adc0_dac_val[8] adc0_dac_val[7] adc0_dac_val[6]
+ adc0_dac_val[5] adc0_dac_val[4] adc0_dac_val[3] adc0_dac_val[2] adc0_dac_val[1]
+ adc0_dac_val[0] audiodac_outb_to_analog0[0] audiodac_out_to_analog1[0] porb_h[0]
Xsky130_ef_ip__scomp3v_0 adc1_comp_out vdda0 sky130_ef_ip__scomp3v_0/VINP left_vref
+ adc1_ena vccd0 w_175560_31974# vssa0 w_178222_28294# vssd0 sky130_ef_ip__scomp3v
Xsky130_td_ip__opamp_hp_narrow_2 vdda0 right_hgbw_opamp_out right_hgbw_opamp_ibias
+ right_hgbw_opamp_in_n right_hgbw_opamp_in_p vssa0 vccd0 vssd0 right_hgbw_opamp_ena
+ sky130_td_ip__opamp_hp_narrow
Xsky130_pa_ip__instramp_1 right_instramp_G2[4] right_instramp_G2[3] right_instramp_G2[2]
+ right_instramp_G2[1] right_instramp_G2[0] right_instramp_G1[4] right_instramp_G1[3]
+ right_instramp_G1[2] right_instramp_G1[1] right_instramp_G1[0] right_vref ibias_instr2
+ right_instramp_in_p vccd0 right_instramp_out right_instramp_in_n w_533800_87810#
+ w_533800_84326# w_524052_102828# w_524052_88784# w_543520_84326# w_533772_102830#
+ w_533800_88792# w_524052_103810# w_524052_99332# w_543520_88792# w_543520_102832#
+ w_524052_87802# w_524052_84318# w_533772_103812# w_543520_103814# w_543520_99336#
+ w_533772_99334# w_543520_87810# vdda0 vssa0 vssd0 sky130_pa_ip__instramp
Xsky130_ef_ip__scomp3v_1 adc0_comp_out vdda0 sky130_ef_ip__scomp3v_1/VINP right_vref
+ adc0_ena vccd0 w_232980_32142# vssa0 w_235642_28462# vssd0 sky130_ef_ip__scomp3v
Xsky130_td_ip__opamp_hp_narrow_3 vdda0 right_lp_opamp_out right_lp_opamp_ibias right_lp_opamp_in_n
+ right_lp_opamp_in_p vssa0 vccd0 vssd0 right_lp_opamp_ena sky130_td_ip__opamp_hp_narrow
Xsimple_switch_array_53_0 right_hgbw_opamp_p_to_left_vref left_instramp_n_to_right_vref
+ adc0_to_vbgtc right_hgbw_opamp_p_to_voutref vdda0 vccd0 right_hgbw_opamp_n_to_vinref
+ vccd0 adc1_to_right_vref adc1_to_vbgsc vdda0 right_lp_opamp_n_to_vbgtc left_instramp_n_to_vinref
+ vdda0 vccd0 vdda0 right_hgbw_opamp_n_to_right_vref vccd0 vdda0 ulpcomp_p_to_left_vref
+ comp_p_to_tempsense vccd0 vccd0 left_hgbw_opamp_p_to_tempsense vccd0 adc1_to_vinref
+ vccd0 right_hgbw_opamp_n_to_vbgsc vdda0 vdda0 right_hgbw_opamp_in_n vdda0 ulpcomp_p_to_voutref
+ vccd0 right_lp_opamp_p_to_left_vref left_hgbw_opamp_n_to_right_vref comp_p_to_vbgtc
+ right_hgbw_opamp_in_p vccd0 vccd0 right_lp_opamp_p_to_voutref vccd0 vdda0 vccd0
+ vdda0 right_lp_opamp_n_to_vinref comp_n_to_vbgsc comp_n_to_right_vref vccd0 vdda0
+ left_hgbw_opamp_n_to_vinref right_lp_opamp_n_to_right_vref left_hgbw_opamp_in_p
+ vccd0 vssa0 vdda0 vccd0 left_instramp_p_to_left_vref ulpcomp_p_to_tempsense vccd0
+ vccd0 left_lp_opamp_in_p right_lp_opamp_p_to_tempsense vccd0 vdda0 comp_n_to_vinref
+ vssa0 right_instramp_in_p adc0_to_left_vref vbgtc right_instramp_in_n left_instramp_p_to_voutref
+ vccd0 vdda0 vdda0 vssa0 ulpcomp_p vdda0 vssa0 left_lp_opamp_p_to_left_vref ulpcomp_p_to_vbgtc
+ left_hgbw_opamp_in_n left_lp_opamp_p_to_voutref adc0_to_voutref vssa0 left_lp_opamp_n_to_vinref
+ left_lp_opamp_in_n right_instramp_p_to_left_vref vccd0 ulpcomp_n_to_right_vref ulpcomp_n_to_vbgsc
+ vssa0 vccd0 vssa0 vdda0 right_instramp_p_to_voutref vdda0 vccd0 vdda0 vccd0 voutref
+ vssa0 vdda0 vccd0 vssa0 vdda0 left_lp_opamp_n_to_right_vref ulpcomp_n right_instramp_n_to_vinref
+ left_hgbw_opamp_p_to_left_vref vdda0 right_instramp_p_to_tempsense vccd0 vccd0 vssa0
+ left_hgbw_opamp_n_to_vbgtc ulpcomp_n_to_vinref vssa0 vinref vssa0 comp_p vssa0 vssa0
+ vbgsc vdda0 right_instramp_n_to_right_vref adc0 vssa0 vssa0 vssa0 vssa0 vdda0 left_instramp_in_n
+ comp_p_to_left_vref vdda0 adc0_to_tempsense vdda0 right_vref left_instramp_p_to_tempsense
+ right_lp_opamp_in_p vccd0 left_hgbw_opamp_p_to_voutref left_vref vssa0 left_instramp_in_p
+ left_lp_opamp_n_to_vbgsc vssa0 vccd0 vdda0 adc1 right_lp_opamp_in_n vssa0 tempsense_out
+ vssa0 vssa0 vssa0 vdda0 vssa0 vdda0 vssa0 vssa0 vssa0 vdda0 comp_p_to_voutref vssa0
+ comp_n vssa0 vccd0 vssd0 simple_switch_array_53
Xsimple_switch_array_16_0 vdda0 left_instramp_n_to_sio1 left_lp_opamp_in_p comp_p
+ right_lp_opamp_p_to_sio0 left_lp_opamp_in_n left_lp_opamp_n_to_sio1 comp_n comp_n_to_sio1
+ left_lp_opamp_p_to_sio0 left_hgbw_opamp_p_to_sio0 right_hgbw_opamp_n_to_sio1 right_lp_opamp_n_to_sio1
+ right_hgbw_opamp_in_p right_instramp_n_to_sio1 right_hgbw_opamp_in_n left_hgbw_opamp_in_p
+ left_hgbw_opamp_in_n right_instramp_p_to_sio0 ulpcomp_p_to_sio0 right_instramp_in_p
+ left_instramp_p_to_sio0 right_instramp_in_n ulpcomp_p right_hgbw_opamp_p_to_sio0
+ ulpcomp_n sio1_core right_lp_opamp_in_p sio0_core left_hgbw_opamp_n_to_sio1 left_instramp_in_p
+ right_lp_opamp_in_n vccd0 comp_p_to_sio0 left_instramp_in_n ulpcomp_n_to_sio1 vssa0
+ vssd0 simple_switch_array_16
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_0[0] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_0[1] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_0[2] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_0[3] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_0[4] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_0[5] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_0[6] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_0[7] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_0[8] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_0[9] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[0|0] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[1|0] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[2|0] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[3|0] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[4|0] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[5|0] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[0|1] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[1|1] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[2|1] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[3|1] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[4|1] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[5|1] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[0|2] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[1|2] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[2|2] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[3|2] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[4|2] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_1[5|2] vssio vbgpwr sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_ef_ip__idac3v_8bit_0 idac_value[6] idac_value[3] idac_value[2] idac_value[0]
+ idac_value[1] idac_value[5] idac_value[4] idac_value[7] ibias_ref_select idac_ena
+ vbg idac_src vdda1 vdda0 idac_snk vccd0 vssd0 vssa0 sky130_ef_ip__idac3v_8bit
Xsky130_fd_io__top_pwrdetv2_0 vssa1 vssa1 sky130_fd_io__top_pwrdetv2_0/out3_vddio_hv
+ sky130_fd_io__top_pwrdetv2_0/out1_vddio_hv sky130_fd_io__top_pwrdetv2_0/out2_vddio_hv
+ sky130_fd_io__top_pwrdetv2_0/out2_vddd_hv sky130_fd_io__top_pwrdetv2_0/out1_vddd_hv
+ vssa1 vccd1_pwr_good vdda1_pwr_good sky130_fd_io__top_pwrdetv2_0/tie_lo_esd porb_h[0]
+ sky130_fd_io__top_pwrdetv2_0/out3_vddd_hv vssa1 vssa1 vssa1 vssd1 vccd0 vccd0 vssa1
+ vccd1 vdda1 vssd0 sky130_fd_io__top_pwrdetv2
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[0] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[1] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[2] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[3] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[4] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[5] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[6] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[7] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[8] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[9] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[10] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[11] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[12] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[13] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[14] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_2[15] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_io__top_pwrdetv2_1 vssa2 vssa2 sky130_fd_io__top_pwrdetv2_1/out3_vddio_hv
+ sky130_fd_io__top_pwrdetv2_1/out1_vddio_hv sky130_fd_io__top_pwrdetv2_1/out2_vddio_hv
+ sky130_fd_io__top_pwrdetv2_1/out2_vddd_hv sky130_fd_io__top_pwrdetv2_1/out1_vddd_hv
+ vssa2 vccd2_pwr_good vdda2_pwr_good sky130_fd_io__top_pwrdetv2_1/tie_lo_esd porb_h[0]
+ sky130_fd_io__top_pwrdetv2_1/out3_vddd_hv vssa2 vssa2 vssa2 vssd2 vccd0 vccd0 vssa2
+ vccd2 vdda2 vssd0 sky130_fd_io__top_pwrdetv2
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_3[0] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_3[1] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_3[2] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_3[3] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_3[4] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_3[5] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_3[6] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_3[7] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_3[8] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_3[9] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_ajc_ip__brownout_0 vdda0 sky130_ajc_ip__brownout_0/outb vccd0 sky130_ajc_ip__brownout_0/osc_ck
+ brownout_unfilt vbg brownout_otrip[2] brownout_otrip[1] brownout_otrip[0] sky130_ajc_ip__brownout_0/itest
+ brownout_filt brownout_vtrip[2] brownout_vtrip[1] brownout_vtrip[0] sky130_ajc_ip__brownout_0/vin_brout
+ brownout_ena brownout_rc_ena sky130_ajc_ip__brownout_0/vin_vunder brownout_rc_dis
+ brownout_timeout brownout_vunder brownout_oneshot brownout_isrc_sel brownout_ibias
+ sky130_ajc_ip__brownout_0/brownout_ana_0/comparator_1/vt sky130_ajc_ip__brownout_0/brownout_ana_0/comparator_0/vt
+ vssa0 vssd0 sky130_ajc_ip__brownout
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[0] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[1] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[2] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[3] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[4] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[5] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[6] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[7] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[8] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[9] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[10] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[11] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[12] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[13] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_4[14] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_5[0] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_5[1] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_5[2] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_5[3] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_5[4] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_5[5] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_5[6] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_5[7] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_5[8] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_5[9] vdda0 vssa0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_6[0] vssd0 vccd0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_6[1] vssd0 vccd0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_6[2] vssd0 vccd0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_6[3] vssd0 vccd0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_6[4] vssd0 vccd0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_6[5] vssd0 vccd0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_6[6] vssd0 vccd0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_6[7] vssd0 vccd0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_6[8] vssd0 vccd0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_6[9] vssd0 vccd0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_7[0] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_7[1] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_7[2] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_7[3] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_7[4] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_7[5] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_7[6] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_7[7] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_7[8] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_7[9] vssa0 vdda0 sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_am_ip__ldo_01v8_0 vddio vbgpwr vssio ldo_ena vbg ldo_ref_sel vccd0 vssd0 sky130_am_ip__ldo_01v8
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[0] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[1] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[2] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[3] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[4] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[5] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[6] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[7] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[8] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[9] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[10] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[11] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[12] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[13] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[14] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_8[15] vssio vddio sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_9[0|0] vssio vcmosref sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_9[1|0] vssio vcmosref sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_9[2|0] vssio vcmosref sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_9[3|0] vssio vcmosref sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_9[4|0] vssio vcmosref sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_9[0|1] vssio vcmosref sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_9[1|1] vssio vcmosref sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_9[2|1] vssio vcmosref sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_9[3|1] vssio vcmosref sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsky130_fd_pr__cap_mim_m3_2_KB5CJD_9[4|1] vssio vcmosref sky130_fd_pr__cap_mim_m3_2_KB5CJD
Xsimple_switch_array_3_0 right_instramp_in_p left_lp_opamp_n_to_rheostat_tap left_lp_opamp_in_n
+ right_instramp_n_to_left_rheostat2_out sky130_ef_ip__rheostat_8bit_4/Vhigh right_instramp_p_to_left_rheostat2_out
+ right_instramp_in_n vssa0 sky130_ef_ip__rheostat_8bit_4/out sky130_ef_ip__rheostat_8bit_4/Vhigh
+ vccd0 vdda0 vssd0 simple_switch_array_3
Xsimple_switch_array_3_1 left_hgbw_opamp_in_n left_instramp_p_to_left_rheostat1_out
+ left_instramp_in_p left_instramp_n_to_left_rheostat1_out sky130_ef_ip__rheostat_8bit_0/Vhigh
+ left_hgbw_opamp_n_to_rheostat_tap left_instramp_in_n vssa0 sky130_ef_ip__rheostat_8bit_0/Vhigh
+ sky130_ef_ip__rheostat_8bit_0/out vccd0 vdda0 vssd0 simple_switch_array_3
Xsimple_switch_array_3_2 right_instramp_in_p right_hgbw_opamp_n_to_rheostat_tap right_hgbw_opamp_in_n
+ right_instramp_n_to_right_rheostat1_out sky130_ef_ip__rheostat_8bit_3/Vhigh right_instramp_p_to_right_rheostat1_out
+ right_instramp_in_n vssa0 sky130_ef_ip__rheostat_8bit_3/out sky130_ef_ip__rheostat_8bit_3/Vhigh
+ vccd0 vdda0 vssd0 simple_switch_array_3
Xsky130_ak_ip__cmos_vref_0 vcmosref vbgpwr bandgap_ena vbgsc vbgtc bandgap_trim[3]
+ bandgap_trim[2] bandgap_trim[1] bandgap_trim[0] sky130_ak_ip__cmos_vref_0/vptat
+ vccd0 vssd0 vssio sky130_ak_ip__cmos_vref
Xsky130_sw_ip__por_0 por vddio vccd0 porb vssd0 porb_h[0] porb_h[1] vssio sky130_sw_ip__por
Xsimple_switch_array_3_3 right_lp_opamp_in_n left_instramp_p_to_right_rheostat2_out
+ left_instramp_in_p left_instramp_n_to_right_rheostat2_out sky130_ef_ip__rheostat_8bit_2/Vhigh
+ right_lp_opamp_n_to_rheostat_tap left_instramp_in_n vssa0 sky130_ef_ip__rheostat_8bit_2/Vhigh
+ sky130_ef_ip__rheostat_8bit_2/out vccd0 vdda0 vssd0 simple_switch_array_3
Xswitch_array_18_0 left_lp_opamp_to_comp_n[0] right_instramp_out right_instramp_to_comp_n[1]
+ left_instramp_out left_hgbw_opamp_to_adc0[0] right_lp_opamp_to_adc0[0] right_hgbw_opamp_out
+ right_instramp_to_adc1[0] right_hgbw_opamp_to_adc1[1] vccd0 vssd0 right_lp_opamp_to_comp_p[1]
+ left_instramp_to_comp_p[0] left_lp_opamp_to_ulpcomp_n[0] vdda0 left_lp_opamp_to_comp_n[1]
+ left_instramp_to_adc0[0] right_lp_opamp_to_adc0[1] left_hgbw_opamp_to_ulpcomp_p[1]
+ left_instramp_to_ulpcomp_p[0] left_hgbw_opamp_out left_hgbw_opamp_to_ulpcomp_p[0]
+ right_hgbw_opamp_to_ulpcomp_n[1] right_hgbw_opamp_to_ulpcomp_n[0] comp_p right_hgbw_opamp_to_adc1[0]
+ adc0 left_lp_opamp_to_ulpcomp_n[1] right_hgbw_opamp_to_comp_n[1] right_lp_opamp_to_comp_p[0]
+ left_hgbw_opamp_to_comp_p[0] left_hgbw_opamp_to_comp_p[1] left_lp_opamp_to_adc1[1]
+ right_lp_opamp_to_ulpcomp_p[0] left_hgbw_opamp_to_adc0[1] comp_n left_instramp_to_ulpcomp_p[1]
+ ulpcomp_p right_instramp_to_ulpcomp_n[1] adc1 right_lp_opamp_to_ulpcomp_p[1] left_instramp_to_adc0[1]
+ ulpcomp_n left_lp_opamp_to_adc1[0] right_lp_opamp_out right_instramp_to_adc1[1]
+ right_hgbw_opamp_to_comp_n[0] left_instramp_to_comp_p[1] right_instramp_to_comp_n[0]
+ left_lp_opamp_out right_instramp_to_ulpcomp_n[0] vssa0 switch_array_18
Xsky130_iic_ip__audiodac_drv_lite_0 audiodac_in audiodac_inb audiodac_out audiodac_outb
+ vccd0 vdda0 vssa0 sky130_iic_ip__audiodac_drv_lite
Xsky130_vbl_ip__overvoltage_0 vdda0 vccd0 overvoltage_ena overvoltage_trim[3] ibias_ov
+ overvoltage_trim[2] overvoltage_out vbg overvoltage_trim[1] overvoltage_trim[0]
+ vssd0 vssa0 sky130_vbl_ip__overvoltage
Xswitch_array_4_10 left_lp_opamp_n_to_gpio5_5[1] left_lp_opamp_n_to_gpio5_5[0] left_lp_opamp_p_to_gpio5_4[1]
+ left_lp_opamp_p_to_gpio5_4[0] left_instramp_p_to_gpio5_6[1] left_instramp_p_to_gpio5_6[0]
+ left_instramp_n_to_gpio5_7[1] left_instramp_n_to_gpio5_7[0] left_lp_opamp_in_n gpio5_5
+ gpio5_4 left_instramp_in_p gpio5_6 left_instramp_in_n gpio5_7 vssd0 vdda0 vccd0
+ left_lp_opamp_in_p vssa0 switch_array_4
Xswitch_array_4_11 ulpcomp_n_to_gpio6_1[1] ulpcomp_n_to_gpio6_1[0] ulpcomp_p_to_gpio6_0[1]
+ ulpcomp_p_to_gpio6_0[0] comp_p_to_gpio6_2[1] comp_p_to_gpio6_2[0] comp_n_to_gpio6_3[1]
+ comp_n_to_gpio6_3[0] ulpcomp_n gpio6_1 gpio6_0 comp_p gpio6_2 comp_n gpio6_3 vssd0
+ vdda0 vccd0 ulpcomp_p vssa0 switch_array_4
Xsimple_switch_array_15_0 user_vinref vdda0 vbgtc_to_user comp_p vbgsc_to_user user_to_adc1[1]
+ vinref_to_user right_vref_to_user comp_n left_vref user_to_ulpcomp_n[1] user_to_comp_n[0]
+ dac0_to_user right_vref user_adc1 user_vbgsc dac1 user_adc0 user_vbgtc user_to_ulpcomp_p[0]
+ dac0 vinref dac1_to_user tempsense_out user_to_adc0[1] user_tempsense vbgsc vbgtc
+ user_to_adc1[0] user_to_comp_p[1] voutref_to_user user_to_ulpcomp_n[0] user_dac1
+ user_dac0 left_vref_to_user ulpcomp_p user_left_vref tempsense_to_user ulpcomp_n
+ user_to_adc0[0] user_to_comp_n[1] user_comp_p user_right_vref user_ulpcomp_p user_comp_n
+ user_to_comp_p[0] user_to_ulpcomp_p[1] user_ulpcomp_n adc1 adc0 vccd0 voutref vssa0
+ vssd0 user_voutref simple_switch_array_15
Xsimple_switch_array_8_0 comp_p ulpcomp_p ulpcomp_p_to_dac0 right_hgbw_opamp_p_to_dac0
+ right_hgbw_opamp_in_n right_lp_opamp_in_n comp_n_to_dac1 right_lp_opamp_n_to_dac1
+ ulpcomp_n_to_dac1 right_hgbw_opamp_n_to_dac1 right_hgbw_opamp_in_p comp_n right_lp_opamp_p_to_dac0
+ right_lp_opamp_in_p comp_p_to_dac0 vccd0 dac0 ulpcomp_n vssa0 dac1 vdda0 vssd0 simple_switch_array_8
Xsky130_ef_ip__rheostat_8bit_0 left_rheostat1_b[0] left_rheostat1_b[1] left_rheostat1_b[2]
+ left_rheostat1_b[3] left_rheostat1_b[4] left_rheostat1_b[5] left_rheostat1_b[6]
+ left_rheostat1_b[7] sky130_ef_ip__rheostat_8bit_0/out vdda0 vccd0 sky130_ef_ip__rheostat_8bit_0/Vhigh
+ vssa0 left_hgbw_opamp_out vssd0 sky130_ef_ip__rheostat_8bit
Xswitch_array_14_1 vccd0 left_hgbw_opamp_out right_instramp_out left_lp_opamp_to_analog0[1]
+ analog1_connect[0] right_hgbw_opamp_to_analog0[0] left_instramp_out right_hgbw_opamp_out
+ left_hgbw_opamp_to_analog1[0] amuxbus_a_n vdda0 vssd0 left_instramp_to_amuxbusB[0]
+ right_instramp_to_analog0[0] right_hgbw_opamp_to_amuxbusA[0] right_lp_opamp_to_analog1[0]
+ analog1 right_instramp_to_amuxbusA[0] analog0 left_lp_opamp_to_analog0[0] analog1_core
+ left_instramp_to_analog1[0] analog0_core left_instramp_to_analog1[1] amuxbus_b_n
+ analog0_connect[0] left_lp_opamp_to_amuxbusA[0] analog0_connect[1] left_hgbw_opamp_to_amuxbusB[0]
+ right_hgbw_opamp_to_analog0[1] left_lp_opamp_to_amuxbusA[1] analog1_connect[1] left_hgbw_opamp_to_analog1[1]
+ right_lp_opamp_to_amuxbusB[0] left_instramp_to_amuxbusB[1] right_instramp_to_analog0[1]
+ right_instramp_to_amuxbusA[1] right_hgbw_opamp_to_amuxbusA[1] right_lp_opamp_to_analog1[1]
+ left_hgbw_opamp_to_amuxbusB[1] right_lp_opamp_out right_lp_opamp_to_amuxbusB[1]
+ left_lp_opamp_out vssa0 switch_array_14
Xswitch_array_4_0 left_instramp_to_gpio4_4[1] left_instramp_to_gpio4_4[0] left_hgbw_opamp_to_gpio4_5[1]
+ left_hgbw_opamp_to_gpio4_5[0] right_lp_opamp_to_gpio4_7[1] right_lp_opamp_to_gpio4_7[0]
+ right_hgbw_opamp_to_gpio4_6[1] right_hgbw_opamp_to_gpio4_6[0] left_instramp_out
+ gpio4_4 gpio4_5 right_lp_opamp_out gpio4_7 right_hgbw_opamp_out gpio4_6 vssd0 vdda0
+ vccd0 left_hgbw_opamp_out vssa0 switch_array_4
Xswitch_array_4_1 left_lp_opamp_to_gpio4_0[1] left_lp_opamp_to_gpio4_0[0] left_hgbw_opamp_to_gpio4_1[1]
+ left_hgbw_opamp_to_gpio4_1[0] right_lp_opamp_to_gpio4_3[1] right_lp_opamp_to_gpio4_3[0]
+ right_hgbw_opamp_to_gpio4_2[1] right_hgbw_opamp_to_gpio4_2[0] left_lp_opamp_out
+ gpio4_0 gpio4_1 right_lp_opamp_out gpio4_3 right_hgbw_opamp_out gpio4_2 vssd0 vdda0
+ vccd0 left_hgbw_opamp_out vssa0 switch_array_4
Xsky130_ef_ip__rheostat_8bit_2 right_rheostat2_b[0] right_rheostat2_b[1] right_rheostat2_b[2]
+ right_rheostat2_b[3] right_rheostat2_b[4] right_rheostat2_b[5] right_rheostat2_b[6]
+ right_rheostat2_b[7] sky130_ef_ip__rheostat_8bit_2/out vdda0 vccd0 sky130_ef_ip__rheostat_8bit_2/Vhigh
+ vssa0 right_lp_opamp_out vssd0 sky130_ef_ip__rheostat_8bit
Xswitch_array_4_2 left_lp_opamp_to_gpio3_4[1] left_lp_opamp_to_gpio3_4[0] left_hgbw_opamp_to_gpio3_5[1]
+ left_hgbw_opamp_to_gpio3_5[0] right_lp_opamp_to_gpio3_7[1] right_lp_opamp_to_gpio3_7[0]
+ right_hgbw_opamp_to_gpio3_6[1] right_hgbw_opamp_to_gpio3_6[0] left_lp_opamp_out
+ gpio3_4 gpio3_5 right_lp_opamp_out gpio3_7 right_hgbw_opamp_out gpio3_6 vssd0 vdda0
+ vccd0 left_hgbw_opamp_out vssa0 switch_array_4
Xsimple_switch_array_6_0 left_hgbw_opamp_in_p left_lp_opamp_in_n adc1 dac1 adc0_to_dac0
+ left_lp_opamp_p_to_dac0 left_hgbw_opamp_p_to_dac0 left_lp_opamp_n_to_dac1 adc0 vdda0
+ left_lp_opamp_in_p vccd0 dac0 adc1_to_dac1 left_hgbw_opamp_in_n left_hgbw_opamp_n_to_dac1
+ vssa0 vssd0 simple_switch_array_6
Xsky130_ef_ip__rheostat_8bit_3 right_rheostat1_b[0] right_rheostat1_b[1] right_rheostat1_b[2]
+ right_rheostat1_b[3] right_rheostat1_b[4] right_rheostat1_b[5] right_rheostat1_b[6]
+ right_rheostat1_b[7] sky130_ef_ip__rheostat_8bit_3/out vdda0 vccd0 sky130_ef_ip__rheostat_8bit_3/Vhigh
+ vssa0 right_hgbw_opamp_out vssd0 sky130_ef_ip__rheostat_8bit
Xsky130_od_ip__tempsensor_ext_vp_0 simple_analog_mux_sel1v8_0/inB simple_analog_mux_sel1v8_0/inA
+ tempsense_ena vbg vccd0 vssd0 sky130_od_ip__tempsensor_ext_vp
Xswitch_array_4_3 right_lp_opamp_to_gpio3_3[1] right_lp_opamp_to_gpio3_3[0] right_hgbw_opamp_to_gpio3_2[1]
+ right_hgbw_opamp_to_gpio3_2[0] right_instramp_to_gpio3_0[1] right_instramp_to_gpio3_0[0]
+ left_hgbw_opamp_to_gpio3_1[1] left_hgbw_opamp_to_gpio3_1[0] right_lp_opamp_out gpio3_3
+ gpio3_2 right_instramp_out gpio3_0 left_hgbw_opamp_out gpio3_1 vssd0 vdda0 vccd0
+ right_hgbw_opamp_out vssa0 switch_array_4
Xswitch_array_2_0 audiodac_out_to_analog1[1] audiodac_out_to_analog1[0] audiodac_outb_to_analog0[1]
+ audiodac_outb_to_analog0[0] audiodac_out audiodac_outb analog0_core vdda0 vssd0
+ analog1_core vccd0 vssa0 switch_array_2
Xsky130_ef_ip__rheostat_8bit_4 left_rheostat2_b[0] left_rheostat2_b[1] left_rheostat2_b[2]
+ left_rheostat2_b[3] left_rheostat2_b[4] left_rheostat2_b[5] left_rheostat2_b[6]
+ left_rheostat2_b[7] sky130_ef_ip__rheostat_8bit_4/out vdda0 vccd0 sky130_ef_ip__rheostat_8bit_4/Vhigh
+ vssa0 left_lp_opamp_out vssd0 sky130_ef_ip__rheostat_8bit
Xswitch_array_4_4 right_hgbw_opamp_n_to_gpio2_2[1] right_hgbw_opamp_n_to_gpio2_2[0]
+ right_hgbw_opamp_p_to_gpio2_3[1] right_hgbw_opamp_p_to_gpio2_3[0] dac_refl_to_gpio1_0[1]
+ dac_refl_to_gpio1_0[0] dac_refh_to_gpio1_1[1] dac_refh_to_gpio1_1[0] right_hgbw_opamp_in_n
+ gpio2_2 gpio2_3 dac_vrefL gpio1_0 dac_vrefH gpio1_1 vssd0 vdda0 vccd0 right_hgbw_opamp_in_p
+ vssa0 switch_array_4
Xswitch_array_2_1 ibias_test_to_gpio1_2[1] ibias_test_to_gpio1_2[0] vbg_test_to_gpio1_1[1]
+ vbg_test_to_gpio1_1[0] ibias_test vbg gpio1_1 vdda0 vssd0 gpio1_2 vccd0 vssa0 switch_array_2
Xsimple_analog_mux_sel1v8_0 simple_analog_mux_sel1v8_0/inA tempsense_out vdda0 vccd0
+ tempsense_sel simple_analog_mux_sel1v8_0/inB vssd0 vssa0 simple_analog_mux_sel1v8
Xswitch_array_4_5 ulpcomp_n_to_gpio1_6[1] ulpcomp_n_to_gpio1_6[0] ulpcomp_p_to_gpio1_7[1]
+ ulpcomp_p_to_gpio1_7[0] left_hgbw_opamp_n_to_gpio2_0[1] left_hgbw_opamp_n_to_gpio2_0[0]
+ left_hgbw_opamp_p_to_gpio2_1[1] left_hgbw_opamp_p_to_gpio2_1[0] ulpcomp_n gpio1_6
+ gpio1_7 left_hgbw_opamp_in_n gpio2_0 left_hgbw_opamp_in_p gpio2_1 vssd0 vdda0 vccd0
+ ulpcomp_p vssa0 switch_array_4
Xswitch_array_2_2 idac_to_gpio1_3[1] idac_to_gpio1_3[0] idac_to_gpio1_2[1] idac_to_gpio1_2[0]
+ idac_snk idac_src gpio1_2 vdda0 vssd0 gpio1_3 vccd0 vssa0 switch_array_2
Xsimple_analog_mux_sel1v8_1 simple_analog_mux_sel1v8_1/inA vbg vdda0 vccd0 bandgap_sel
+ vcmosref vssd0 vssa0 simple_analog_mux_sel1v8
Xswitch_array_4_6 right_hgbw_opamp_n_to_gpio5_1[1] right_hgbw_opamp_n_to_gpio5_1[0]
+ right_hgbw_opamp_p_to_gpio5_0[1] right_hgbw_opamp_p_to_gpio5_0[0] left_hgbw_opamp_p_to_gpio5_2[1]
+ left_hgbw_opamp_p_to_gpio5_2[0] left_hgbw_opamp_n_to_gpio5_3[1] left_hgbw_opamp_n_to_gpio5_3[0]
+ right_hgbw_opamp_in_n gpio5_1 gpio5_0 left_hgbw_opamp_in_p gpio5_2 left_hgbw_opamp_in_n
+ gpio5_3 vssd0 vdda0 vccd0 right_hgbw_opamp_in_p vssa0 switch_array_4
Xswitch_array_2_3 sio1_connect[1] sio1_connect[0] sio0_connect[1] sio0_connect[0]
+ sio1_core sio0_core sio0 vdda0 vssd0 sio1 vccd0 vssa0 switch_array_2
Xsky130_ak_ip__comparator_0 comp_p comp_n vdda0 comp_ena comp_hyst[1] comp_hyst[0]
+ comp_trim[5] comp_trim[4] comp_trim[3] comp_trim[2] comp_trim[1] comp_trim[0] comp_out
+ vccd0 ibias_comp vssd0 vssa0 sky130_ak_ip__comparator
Xsky130_icrg_ip__ulpcomp2_0 vdda0 ulpcomp_ena ulpcomp_out ulpcomp_n ulpcomp_p vssd0
+ ulpcomp_clk vccd0 vssa0 w_364506_55555# sky130_icrg_ip__ulpcomp2
Xswitch_array_4_7 adc1_to_gpio6_5[1] adc1_to_gpio6_5[0] adc0_to_gpio6_4[1] adc0_to_gpio6_4[0]
+ adc_refh_to_gpio6_6[1] adc_refh_to_gpio6_6[0] adc_refl_to_gpio6_7[1] adc_refl_to_gpio6_7[0]
+ adc1 gpio6_5 gpio6_4 adc_vrefH gpio6_6 adc_vrefL gpio6_7 vssd0 vdda0 vccd0 adc0
+ vssa0 switch_array_4
Xswitch_array_4_8 right_instramp_p_to_gpio2_7[1] right_instramp_p_to_gpio2_7[0] right_instramp_n_to_gpio2_6[1]
+ right_instramp_n_to_gpio2_6[0] right_lp_opamp_p_to_gpio2_5[1] right_lp_opamp_p_to_gpio2_5[0]
+ right_lp_opamp_n_to_gpio2_4[1] right_lp_opamp_n_to_gpio2_4[0] right_instramp_in_p
+ gpio2_7 gpio2_6 right_lp_opamp_in_p gpio2_5 right_lp_opamp_in_n gpio2_4 vssd0 vdda0
+ vccd0 right_instramp_in_n vssa0 switch_array_4
Xsky130_ef_ip__cdac3v_12bit_0 adc1_dac_val[2] adc1_dac_val[3] adc1_dac_val[4] adc1_dac_val[5]
+ adc1_dac_val[6] adc1_dac_val[7] adc1_dac_val[8] adc1_dac_val[9] vdda0 vccd0 sky130_ef_ip__scomp3v_0/VINP
+ adc1_reset adc1_dac_val[10] adc1_dac_val[11] sky130_ef_ip__cdac3v_12bit_0/OUTNC
+ adc1_dac_val[0] adc1_dac_val[1] vinref adc1 adc1_hold left_vref adc_vrefL adc_vrefH
+ vssa0 vssd0 sky130_ef_ip__cdac3v_12bit
Xswitch_array_4_9 adc1_to_gpio1_2[1] adc1_to_gpio1_2[0] adc0_to_gpio1_3[1] adc0_to_gpio1_3[0]
+ comp_n_to_gpio1_4[1] comp_n_to_gpio1_4[0] comp_p_to_gpio1_5[1] comp_p_to_gpio1_5[0]
+ adc1 gpio1_2 gpio1_3 comp_n gpio1_4 comp_p gpio1_5 vssd0 vdda0 vccd0 adc0 vssa0
+ switch_array_4
Xsky130_ef_ip__rdac3v_8bit_0 rdac0_value[0] rdac0_value[1] rdac0_value[2] rdac0_value[3]
+ rdac0_value[4] rdac0_value[5] rdac0_value[6] rdac0_value[7] dac0 vdda0 rdac0_ena
+ vccd0 dac_vrefH dac_vrefL vssa0 vssd0 sky130_ef_ip__rdac3v_8bit
Xsky130_ef_ip__cdac3v_12bit_1 adc0_dac_val[2] adc0_dac_val[3] adc0_dac_val[4] adc0_dac_val[5]
+ adc0_dac_val[6] adc0_dac_val[7] adc0_dac_val[8] adc0_dac_val[9] vdda0 vccd0 sky130_ef_ip__scomp3v_1/VINP
+ adc0_reset adc0_dac_val[10] adc0_dac_val[11] sky130_ef_ip__cdac3v_12bit_1/OUTNC
+ adc0_dac_val[0] adc0_dac_val[1] voutref adc0 adc0_hold right_vref adc_vrefL adc_vrefH
+ vssa0 vssd0 sky130_ef_ip__cdac3v_12bit
Xsimple_switch_array_32_0 vdda0 left_lp_opamp_in_p right_instramp_p_to_analog0 comp_p
+ left_lp_opamp_in_n left_hgbw_opamp_p_to_analog0 comp_n left_hgbw_opamp_n_to_analog1
+ ulpcomp_p_to_analog1 left_instramp_n_to_analog1 dac1 ulpcomp_n_to_analog0 dac0 amuxbus_b_n
+ amuxbus_a_n right_instramp_n_to_amuxbusB left_lp_opamp_p_to_amuxbusA left_hgbw_opamp_p_to_amuxbusA
+ analog0_core right_hgbw_opamp_in_p adc0_to_analog1 dac1_to_analog0 right_hgbw_opamp_in_n
+ right_lp_opamp_n_to_analog1 left_hgbw_opamp_in_p comp_p_to_analog1 right_lp_opamp_p_to_amuxbusA
+ right_lp_opamp_p_to_analog0 left_hgbw_opamp_in_n left_instramp_n_to_amuxbusB left_lp_opamp_n_to_amuxbusB
+ comp_n_to_analog0 adc1_to_analog0 right_instramp_in_p dac0_to_analog1 left_lp_opamp_n_to_analog1
+ right_instramp_in_n left_instramp_p_to_analog0 left_instramp_p_to_amuxbusA ulpcomp_p
+ right_hgbw_opamp_p_to_analog0 right_lp_opamp_n_to_amuxbusB ulpcomp_n right_hgbw_opamp_n_to_amuxbusB
+ left_hgbw_opamp_n_to_amuxbusB right_lp_opamp_in_p right_hgbw_opamp_n_to_analog1
+ left_instramp_in_p adc1 right_instramp_n_to_analog1 right_lp_opamp_in_n right_hgbw_opamp_p_to_amuxbusA
+ adc0 vccd0 left_lp_opamp_p_to_analog0 left_instramp_in_n right_instramp_p_to_amuxbusA
+ vssa0 analog1_core vssd0 simple_switch_array_32
Xsky130_ef_ip__biasgen4_0 ibias_ena ibias_ref_select vccd0 vdda0 vbg ibias_snk_ena[3]
+ ibias_snk_ena[2] ibias_snk_ena[1] ibias_snk_ena[0] ibias_src_ena[2] ibias_src_ena[1]
+ ibias_src_ena[12] ibias_src_ena[0] ibias_src_ena[5] ibias_src_ena[3] ibias_src_ena[4]
+ ibias_src_ena[10] ibias_src_ena[9] ibias_src_ena[7] ibias_src_ena[8] ibias_src_ena[17]
+ ibias_src_ena[16] ibias_src_ena[11] ibias_src_ena[15] ibias_src_ena[23] ibias_src_ena[22]
+ ibias_src_ena[20] ibias_src_ena[21] ibias_src_ena[18] ibias_src_ena[14] ibias_src_ena[19]
+ ibias_src_ena[13] ibias_src_ena[6] ibias_lsxo left_lp_opamp_ibias right_lp_opamp_ibias
+ left_hgbw_opamp_ibias right_hgbw_opamp_ibias ibias_instr1 ibias_instr2 ibias_ov
+ user_ibias50 ibias_test brownout_ibias ibias_hsxo ibias_idac vdda1 ibias_comp sky130_cw_ip__bandgap_nobias_0/bias
+ user_ibias100 vssd0 vssa0 sky130_ef_ip__biasgen4
Xsky130_ef_ip__rdac3v_8bit_1 rdac1_value[0] rdac1_value[1] rdac1_value[2] rdac1_value[3]
+ rdac1_value[4] rdac1_value[5] rdac1_value[6] rdac1_value[7] dac1 vdda0 rdac1_ena
+ vccd0 dac_vrefH dac_vrefL vssa0 vssd0 sky130_ef_ip__rdac3v_8bit
Xsky130_cw_ip__bandgap_nobias_0 bandgap_trim[0] bandgap_trim[4] bandgap_trim[6] bandgap_trim[10]
+ bandgap_trim[12] bandgap_trim[14] bandgap_trim[15] bandgap_trim[13] bandgap_trim[11]
+ bandgap_trim[7] bandgap_trim[5] bandgap_trim[3] bandgap_trim[1] bandgap_trim[2]
+ vssd0 sky130_cw_ip__bandgap_nobias_0/bias simple_analog_mux_sel1v8_1/inA bandgap_trim[9]
+ bandgap_trim[8] vccd0 vssd0 sky130_cw_ip__bandgap_nobias
Xsky130_td_ip__opamp_hp_narrow_0 vdda0 left_hgbw_opamp_out left_hgbw_opamp_ibias left_hgbw_opamp_in_n
+ left_hgbw_opamp_in_p vssa0 vccd0 vssd0 left_hgbw_opamp_ena sky130_td_ip__opamp_hp_narrow
Xsky130_td_ip__opamp_hp_narrow_1 vdda0 left_lp_opamp_out left_lp_opamp_ibias left_lp_opamp_in_n
+ left_lp_opamp_in_p vssa0 vccd0 vssd0 left_lp_opamp_ena sky130_td_ip__opamp_hp_narrow
Xsky130_pa_ip__instramp_0 left_instramp_G2[4] left_instramp_G2[3] left_instramp_G2[2]
+ left_instramp_G2[1] left_instramp_G2[0] left_instramp_G1[4] left_instramp_G1[3]
+ left_instramp_G1[2] left_instramp_G1[1] left_instramp_G1[0] left_vref ibias_instr1
+ left_instramp_in_p vccd0 left_instramp_out left_instramp_in_n w_71682_85054# w_71682_81570#
+ w_61934_100072# w_61934_86028# w_81402_81570# w_71654_100074# w_71682_86036# w_61934_101054#
+ w_61934_96576# w_81402_86036# w_81402_100076# w_61934_85046# w_61934_81562# w_71654_101056#
+ w_81402_101058# w_81402_96580# w_71654_96578# w_81402_85054# vdda0 vssa0 vssd0 sky130_pa_ip__instramp
R0 gpio3_4 user_gpio3_4_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R1 gpio4_0 user_gpio4_0_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R2 gpio3_1 user_gpio3_1_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R3 gpio4_6 user_gpio4_6_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R4 gpio3_5 user_gpio3_5_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R5 gpio4_3 user_gpio4_3_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R6 gpio4_1 user_gpio4_1_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R7 gpio3_6 user_gpio3_6_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R8 gpio4_4 user_gpio4_4_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R9 gpio3_2 user_gpio3_2_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R10 gpio4_7 user_gpio4_7_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R11 gpio3_0 user_gpio3_0_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R12 gpio3_7 user_gpio3_7_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R13 gpio4_2 user_gpio4_2_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R14 gpio3_3 user_gpio3_3_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
R15 gpio4_5 user_gpio4_5_analog sky130_fd_pr__res_generic_m4 w=0.64 l=0.23
.ends

