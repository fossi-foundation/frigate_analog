VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_to_gpio_top_right
  CLASS COVER ;
  FOREIGN analog_to_gpio_top_right ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.810 BY 157.940 ;
  OBS
      LAYER met2 ;
        RECT 33.710 153.415 35.280 155.585 ;
      LAYER met3 ;
        RECT 33.560 153.210 35.810 155.585 ;
        RECT 33.700 152.580 35.670 153.210 ;
      LAYER met4 ;
        RECT 0.090 157.240 3.290 157.910 ;
        RECT 0.000 156.310 3.290 157.240 ;
        RECT 0.000 4.745 1.000 156.310 ;
        RECT 33.560 154.540 35.810 154.785 ;
        RECT 3.120 153.830 6.320 154.360 ;
        RECT 3.000 152.760 6.320 153.830 ;
        RECT 32.470 152.940 35.810 154.540 ;
        RECT 0.000 0.745 1.600 4.745 ;
        RECT 3.000 0.000 4.000 152.760 ;
        RECT 33.560 152.410 35.810 152.940 ;
        RECT 6.100 150.250 9.300 150.870 ;
        RECT 6.000 149.270 9.300 150.250 ;
        RECT 6.000 4.745 7.000 149.270 ;
        RECT 5.400 0.745 7.000 4.745 ;
      LAYER met5 ;
        RECT -0.030 157.940 3.410 158.030 ;
        RECT -0.030 156.340 35.800 157.940 ;
        RECT -0.030 156.190 3.410 156.340 ;
        RECT 3.000 154.410 6.440 154.480 ;
        RECT 32.350 154.410 35.790 154.660 ;
        RECT 3.000 152.810 35.810 154.410 ;
        RECT 3.000 152.640 6.440 152.810 ;
        RECT 5.980 150.940 9.420 150.990 ;
        RECT 5.980 149.340 35.800 150.940 ;
        RECT 5.980 149.150 9.420 149.340 ;
        RECT 0.000 0.745 7.005 4.745 ;
  END
END analog_to_gpio_top_right
END LIBRARY

