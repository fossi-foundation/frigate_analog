magic
tech sky130A
magscale 1 2
timestamp 1719174692
<< checkpaint >>
rect 542198 73062 542469 73190
<< metal2 >>
rect 542198 73185 542469 73190
rect 542198 73067 542207 73185
rect 542460 73067 542469 73185
rect 542198 73062 542469 73067
<< via2 >>
rect 542207 73067 542460 73185
<< metal3 >>
rect 542198 73185 542469 73190
rect 542198 73067 542207 73185
rect 542460 73067 542469 73185
rect 542198 73062 542469 73067
<< end >>
