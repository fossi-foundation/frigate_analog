magic
tech sky130A
magscale 1 2
timestamp 1724444186
<< metal1 >>
rect -212 2421 -206 2473
rect -154 2465 -148 2473
rect -154 2429 48 2465
rect -154 2421 -148 2429
rect 4304 2421 4310 2473
rect 4362 2465 4368 2473
rect 4362 2429 4768 2465
rect 4362 2421 4368 2429
rect 8820 2421 8826 2473
rect 8878 2465 8884 2473
rect 8878 2429 9286 2465
rect 8878 2421 8884 2429
rect 13336 2421 13342 2473
rect 13394 2465 13400 2473
rect 13394 2429 13795 2465
rect 13394 2421 13400 2429
rect 23060 2419 23066 2471
rect 23118 2463 23124 2471
rect 23118 2427 23422 2463
rect 23118 2419 23124 2427
rect 27576 2419 27582 2471
rect 27634 2463 27640 2471
rect 27634 2427 28157 2463
rect 27634 2419 27640 2427
rect 32092 2419 32098 2471
rect 32150 2463 32156 2471
rect 32150 2427 32675 2463
rect 32150 2419 32156 2427
rect 36608 2419 36614 2471
rect 36666 2463 36672 2471
rect 36666 2427 37183 2463
rect 36666 2419 36672 2427
rect -1 2013 271 2026
rect -1 1883 13 2013
rect 268 1883 271 2013
rect -1 1872 271 1883
rect 4515 2013 4787 2026
rect 4515 1883 4529 2013
rect 4784 1883 4787 2013
rect 4515 1872 4787 1883
rect 9031 2013 9302 2026
rect 9031 1883 9045 2013
rect 9300 1883 9302 2013
rect 9031 1872 9302 1883
rect 13547 2013 13819 2026
rect 13547 1883 13561 2013
rect 13816 1883 13819 2013
rect 13547 1872 13819 1883
rect 23400 2009 23671 2022
rect 23400 1879 23414 2009
rect 23669 1879 23671 2009
rect 23400 1868 23671 1879
rect 27916 2009 28186 2022
rect 27916 1879 27930 2009
rect 28185 1879 28186 2009
rect 27916 1868 28186 1879
rect 32432 2009 32703 2022
rect 32432 1879 32446 2009
rect 32701 1879 32703 2009
rect 32432 1868 32703 1879
rect 36948 2009 37218 2022
rect 36948 1879 36962 2009
rect 37217 1879 37218 2009
rect 36948 1868 37218 1879
<< via1 >>
rect -206 2421 -154 2473
rect 2651 2460 3132 2556
rect 4310 2421 4362 2473
rect 7167 2460 7648 2556
rect 8826 2421 8878 2473
rect 11683 2460 12164 2556
rect 13342 2421 13394 2473
rect 16199 2460 16680 2556
rect 23066 2419 23118 2471
rect 26052 2456 26533 2552
rect 27582 2419 27634 2471
rect 30568 2456 31049 2552
rect 32098 2419 32150 2471
rect 35084 2456 35565 2552
rect 36614 2419 36666 2471
rect 39600 2456 40081 2552
rect 13 1883 268 2013
rect 4529 1883 4784 2013
rect 9045 1883 9300 2013
rect 13561 1883 13816 2013
rect 23414 1879 23669 2009
rect 27930 1879 28185 2009
rect 32446 1879 32701 2009
rect 36962 1879 37217 2009
<< metal2 >>
rect 13996 4537 17036 4541
rect -974 4119 17036 4537
rect 22176 4123 40428 4551
rect -974 4115 13996 4119
rect -974 871 -636 4115
rect 3476 3559 3996 3991
rect 7992 3559 8512 3991
rect 12508 3559 13028 3991
rect 17024 3559 17544 3991
rect 2638 2602 3139 2616
rect 2638 2556 2656 2602
rect 3117 2572 3139 2602
rect 3117 2556 3141 2572
rect -206 2473 -154 2479
rect 2638 2460 2651 2556
rect 3132 2460 3141 2556
rect 2638 2454 2656 2460
rect 3117 2454 3141 2460
rect 2638 2450 3141 2454
rect 2638 2442 3139 2450
rect -206 2415 -154 2421
rect -198 857 -162 2415
rect -1 2013 288 2026
rect -1 1883 13 2013
rect 268 1883 288 2013
rect -1 1872 288 1883
rect 3686 881 3996 3559
rect 7154 2602 7655 2616
rect 7154 2556 7172 2602
rect 7633 2572 7655 2602
rect 7633 2556 7657 2572
rect 4310 2473 4362 2479
rect 7154 2460 7167 2556
rect 7648 2460 7657 2556
rect 7154 2454 7172 2460
rect 7633 2454 7657 2460
rect 7154 2450 7657 2454
rect 7154 2442 7655 2450
rect 4310 2415 4362 2421
rect 4318 857 4354 2415
rect 4515 2013 4804 2026
rect 4515 1883 4529 2013
rect 4784 1883 4804 2013
rect 4515 1872 4804 1883
rect 8202 881 8512 3559
rect 11670 2602 12171 2616
rect 11670 2556 11688 2602
rect 12149 2572 12171 2602
rect 12149 2556 12173 2572
rect 8826 2473 8878 2479
rect 11670 2460 11683 2556
rect 12164 2460 12173 2556
rect 11670 2454 11688 2460
rect 12149 2454 12173 2460
rect 11670 2450 12173 2454
rect 11670 2442 12171 2450
rect 8826 2415 8878 2421
rect 8834 857 8870 2415
rect 9031 2013 9320 2026
rect 9031 1883 9045 2013
rect 9300 1883 9320 2013
rect 9031 1872 9320 1883
rect 12718 881 13028 3559
rect 16186 2602 16687 2616
rect 16186 2556 16204 2602
rect 16665 2572 16687 2602
rect 16665 2556 16689 2572
rect 13342 2473 13394 2479
rect 16186 2460 16199 2556
rect 16680 2460 16689 2556
rect 16186 2454 16204 2460
rect 16665 2454 16689 2460
rect 16186 2450 16689 2454
rect 16186 2442 16687 2450
rect 13342 2415 13394 2421
rect 13350 857 13386 2415
rect 13547 2013 13836 2026
rect 13547 1883 13561 2013
rect 13816 1883 13836 2013
rect 13547 1872 13836 1883
rect 17234 881 17544 3559
rect 22176 885 22514 4123
rect 26824 3579 27344 3991
rect 26876 3559 27344 3579
rect 31340 3559 31860 3991
rect 35856 3559 36376 3991
rect 40372 3559 40892 3991
rect 26039 2598 26540 2612
rect 26039 2552 26057 2598
rect 26518 2568 26540 2598
rect 26518 2552 26542 2568
rect 23066 2471 23118 2477
rect 26039 2456 26052 2552
rect 26533 2456 26542 2552
rect 26039 2450 26057 2456
rect 26518 2450 26542 2456
rect 26039 2446 26542 2450
rect 26039 2438 26540 2446
rect 23066 2413 23118 2419
rect 23074 865 23110 2413
rect 23400 2009 23689 2022
rect 23400 1879 23414 2009
rect 23669 1879 23689 2009
rect 23400 1868 23689 1879
rect 27034 881 27344 3559
rect 30555 2598 31056 2612
rect 30555 2552 30573 2598
rect 31034 2568 31056 2598
rect 31034 2552 31058 2568
rect 27582 2471 27634 2477
rect 30555 2456 30568 2552
rect 31049 2456 31058 2552
rect 30555 2450 30573 2456
rect 31034 2450 31058 2456
rect 30555 2446 31058 2450
rect 30555 2438 31056 2446
rect 27582 2413 27634 2419
rect 27590 865 27626 2413
rect 27916 2009 28205 2022
rect 27916 1879 27930 2009
rect 28185 1879 28205 2009
rect 27916 1868 28205 1879
rect 31550 881 31860 3559
rect 35071 2598 35572 2612
rect 35071 2552 35089 2598
rect 35550 2568 35572 2598
rect 35550 2552 35574 2568
rect 32098 2471 32150 2477
rect 35071 2456 35084 2552
rect 35565 2456 35574 2552
rect 35071 2450 35089 2456
rect 35550 2450 35574 2456
rect 35071 2446 35574 2450
rect 35071 2438 35572 2446
rect 32098 2413 32150 2419
rect 32106 865 32142 2413
rect 32432 2009 32721 2022
rect 32432 1879 32446 2009
rect 32701 1879 32721 2009
rect 32432 1868 32721 1879
rect 36066 881 36376 3559
rect 39587 2598 40088 2612
rect 39587 2552 39605 2598
rect 40066 2568 40088 2598
rect 40066 2552 40090 2568
rect 36614 2471 36666 2477
rect 39587 2456 39600 2552
rect 40081 2456 40090 2552
rect 39587 2450 39605 2456
rect 40066 2450 40090 2456
rect 39587 2446 40090 2450
rect 39587 2438 40088 2446
rect 36614 2413 36666 2419
rect 36622 865 36658 2413
rect 36948 2009 37237 2022
rect 36948 1879 36962 2009
rect 37217 1879 37237 2009
rect 36948 1868 37237 1879
rect 40582 881 40892 3559
<< via2 >>
rect 617 4718 1632 4862
rect 5133 4718 6148 4862
rect 9649 4718 10664 4862
rect 14165 4718 15180 4862
rect 24018 4714 25033 4858
rect 28534 4714 29549 4858
rect 33050 4714 34065 4858
rect 37566 4714 38581 4858
rect 667 3238 1682 3382
rect 2656 2556 3117 2602
rect 2656 2460 3117 2556
rect 2656 2454 3117 2460
rect 13 1883 268 2013
rect 5183 3238 6198 3382
rect 7172 2556 7633 2602
rect 7172 2460 7633 2556
rect 7172 2454 7633 2460
rect 4529 1883 4784 2013
rect 9699 3238 10714 3382
rect 11688 2556 12149 2602
rect 11688 2460 12149 2556
rect 11688 2454 12149 2460
rect 9045 1883 9300 2013
rect 14215 3238 15230 3382
rect 16204 2556 16665 2602
rect 16204 2460 16665 2556
rect 16204 2454 16665 2460
rect 13561 1883 13816 2013
rect 24068 3234 25083 3378
rect 26057 2552 26518 2598
rect 26057 2456 26518 2552
rect 26057 2450 26518 2456
rect 23414 1879 23669 2009
rect 28584 3234 29599 3378
rect 30573 2552 31034 2598
rect 30573 2456 31034 2552
rect 30573 2450 31034 2456
rect 27930 1879 28185 2009
rect 33100 3234 34115 3378
rect 35089 2552 35550 2598
rect 35089 2456 35550 2552
rect 35089 2450 35550 2456
rect 32446 1879 32701 2009
rect 37616 3234 38631 3378
rect 39605 2552 40066 2598
rect 39605 2456 40066 2552
rect 39605 2450 40066 2456
rect 36962 1879 37217 2009
<< metal3 >>
rect 23393 4879 40446 4880
rect -12 4862 40446 4879
rect -12 4718 617 4862
rect 1632 4718 5133 4862
rect 6148 4718 9649 4862
rect 10664 4718 14165 4862
rect 15180 4858 40446 4862
rect 15180 4718 24018 4858
rect -12 4714 24018 4718
rect 25033 4714 28534 4858
rect 29549 4714 33050 4858
rect 34065 4714 37566 4858
rect 38581 4714 40446 4858
rect -12 4703 40446 4714
rect 23393 4696 40446 4703
rect 23390 3406 40443 3412
rect -7 3382 40443 3406
rect -7 3238 667 3382
rect 1682 3238 5183 3382
rect 6198 3238 9699 3382
rect 10714 3238 14215 3382
rect 15230 3378 40443 3382
rect 15230 3238 24068 3378
rect -7 3234 24068 3238
rect 25083 3234 28584 3378
rect 29599 3234 33100 3378
rect 34115 3234 37616 3378
rect 38631 3234 40443 3378
rect -7 3230 40443 3234
rect 23390 3228 40443 3230
rect 24020 3226 25135 3228
rect 28536 3226 29651 3228
rect 33052 3226 34167 3228
rect 37568 3226 38683 3228
rect 23387 2617 40440 2618
rect 26 2602 40440 2617
rect 26 2454 2656 2602
rect 3117 2454 7172 2602
rect 7633 2454 11688 2602
rect 12149 2454 16204 2602
rect 16665 2598 40440 2602
rect 16665 2454 26057 2598
rect 26 2450 26057 2454
rect 26518 2450 30573 2598
rect 31034 2450 35089 2598
rect 35550 2450 39605 2598
rect 40066 2450 40440 2598
rect 26 2441 40440 2450
rect 23387 2434 40440 2441
rect -7 2013 40433 2037
rect -7 1883 13 2013
rect 268 1883 4529 2013
rect 4784 1883 9045 2013
rect 9300 1883 13561 2013
rect 13816 2009 40433 2013
rect 13816 1883 23414 2009
rect -7 1879 23414 1883
rect 23669 1879 27930 2009
rect 28185 1879 32446 2009
rect 32701 1879 36962 2009
rect 37217 1879 40433 2009
rect -7 1861 40433 1879
rect 23380 1853 40433 1861
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_0 ../ip/sky130_ef_ip__analog_switches/mag
array 0 3 4516 0 0 -4248
timestamp 1724439637
transform 1 0 0 0 -1 4529
box -4 -600 3538 3648
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_1
array 0 3 4516 0 0 -4248
timestamp 1724439637
transform 1 0 23400 0 -1 4529
box -4 -600 3538 3648
<< end >>
