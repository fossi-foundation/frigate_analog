magic
tech sky130A
magscale 1 2
timestamp 1720191374
<< metal1 >>
rect 5834 15257 5891 15285
rect 10660 15257 10717 15285
rect 15486 15257 15543 15285
rect 20312 15257 20369 15285
rect 25138 15257 25195 15285
rect 1008 15244 1131 15257
rect 1008 14871 1017 15244
rect 1120 14871 1131 15244
rect 1008 14859 1131 14871
rect 5834 15244 5957 15257
rect 5834 14871 5843 15244
rect 5946 14871 5957 15244
rect 5834 14859 5957 14871
rect 10660 15244 10783 15257
rect 10660 14871 10669 15244
rect 10772 14871 10783 15244
rect 10660 14859 10783 14871
rect 15486 15244 15609 15257
rect 15486 14871 15495 15244
rect 15598 14871 15609 15244
rect 15486 14859 15609 14871
rect 20312 15244 20435 15257
rect 20312 14871 20321 15244
rect 20424 14871 20435 15244
rect 20312 14859 20435 14871
rect 25138 15244 25261 15257
rect 25138 14871 25147 15244
rect 25250 14871 25261 15244
rect 25138 14859 25261 14871
rect 5834 14843 5891 14859
rect 10660 14843 10717 14859
rect 15486 14843 15543 14859
rect 20312 14843 20369 14859
rect 25138 14843 25195 14859
rect 4844 14665 4850 14684
rect 4860 14665 4899 14684
rect 4844 14657 4899 14665
rect 9670 14665 9676 14684
rect 9686 14665 9725 14684
rect 9670 14657 9725 14665
rect 14496 14665 14502 14684
rect 14512 14665 14551 14684
rect 14496 14657 14551 14665
rect 19322 14665 19328 14684
rect 19338 14665 19377 14684
rect 19322 14657 19377 14665
rect 24148 14665 24154 14684
rect 24164 14665 24203 14684
rect 24148 14657 24203 14665
rect -126 14634 64 14657
rect -126 14284 -100 14634
rect 42 14284 64 14634
rect -126 14260 64 14284
rect 4700 14634 4899 14657
rect 4700 14284 4726 14634
rect 4868 14284 4899 14634
rect 4700 14260 4899 14284
rect 9526 14634 9725 14657
rect 9526 14284 9552 14634
rect 9694 14284 9725 14634
rect 9526 14260 9725 14284
rect 14352 14634 14551 14657
rect 14352 14284 14378 14634
rect 14520 14284 14551 14634
rect 14352 14260 14551 14284
rect 19178 14634 19377 14657
rect 19178 14284 19204 14634
rect 19346 14284 19377 14634
rect 19178 14260 19377 14284
rect 24004 14634 24203 14657
rect 24004 14284 24030 14634
rect 24172 14284 24203 14634
rect 24004 14260 24203 14284
rect 4844 14238 4899 14260
rect 9670 14238 9725 14260
rect 14496 14238 14551 14260
rect 19322 14238 19377 14260
rect 24148 14238 24203 14260
rect 1467 10768 1503 11742
rect 1746 10852 1782 11742
rect 4844 11738 5044 11742
rect 5833 11738 6033 11742
rect 6278 10936 6314 11742
rect 6575 11020 6611 11742
rect 9670 11738 9870 11742
rect 10659 11738 10859 11742
rect 11108 11104 11144 11742
rect 11396 11188 11432 11742
rect 14496 11738 14696 11742
rect 15485 11738 15685 11742
rect 15938 11272 15974 11742
rect 16235 11356 16271 11742
rect 19322 11738 19522 11742
rect 20311 11738 20511 11742
rect 20759 11440 20795 11742
rect 21061 11524 21097 11742
rect 24148 11738 24348 11742
rect 25137 11738 25337 11742
rect 25589 11608 25625 11742
rect 25872 11692 25908 11742
rect 25872 11656 28606 11692
rect 25589 11572 28606 11608
rect 21061 11488 28606 11524
rect 20759 11404 28606 11440
rect 16235 11320 28606 11356
rect 15938 11236 28606 11272
rect 11396 11152 28606 11188
rect 11108 11068 28606 11104
rect 6575 10984 28606 11020
rect 6278 10900 28606 10936
rect 1746 10816 28606 10852
rect 1467 10732 28606 10768
rect 1008 9391 1065 9419
rect 5834 9391 5891 9419
rect 10660 9391 10717 9419
rect 15486 9391 15543 9419
rect 20312 9391 20369 9419
rect 25138 9391 25195 9419
rect 1008 9378 1131 9391
rect 1008 9005 1017 9378
rect 1120 9005 1131 9378
rect 1008 8993 1131 9005
rect 5834 9378 5957 9391
rect 5834 9005 5843 9378
rect 5946 9005 5957 9378
rect 5834 8993 5957 9005
rect 10660 9378 10783 9391
rect 10660 9005 10669 9378
rect 10772 9005 10783 9378
rect 10660 8993 10783 9005
rect 15486 9378 15609 9391
rect 15486 9005 15495 9378
rect 15598 9005 15609 9378
rect 15486 8993 15609 9005
rect 20312 9378 20435 9391
rect 20312 9005 20321 9378
rect 20424 9005 20435 9378
rect 20312 8993 20435 9005
rect 25138 9378 25261 9391
rect 25138 9005 25147 9378
rect 25250 9005 25261 9378
rect 25138 8993 25261 9005
rect 1008 8977 1065 8993
rect 5834 8977 5891 8993
rect 10660 8977 10717 8993
rect 15486 8977 15543 8993
rect 20312 8977 20369 8993
rect 25138 8977 25195 8993
rect 18 8799 24 8818
rect 34 8799 73 8818
rect 18 8791 73 8799
rect 4844 8799 4850 8818
rect 4860 8799 4899 8818
rect 4844 8791 4899 8799
rect 9670 8799 9676 8818
rect 9686 8799 9725 8818
rect 9670 8791 9725 8799
rect 14496 8799 14502 8818
rect 14512 8799 14551 8818
rect 14496 8791 14551 8799
rect 19322 8799 19328 8818
rect 19338 8799 19377 8818
rect 19322 8791 19377 8799
rect 24148 8799 24154 8818
rect 24164 8799 24203 8818
rect 24148 8791 24203 8799
rect -126 8768 73 8791
rect -126 8418 -100 8768
rect 42 8418 73 8768
rect -126 8394 73 8418
rect 4700 8768 4899 8791
rect 4700 8418 4726 8768
rect 4868 8418 4899 8768
rect 4700 8394 4899 8418
rect 9526 8768 9725 8791
rect 9526 8418 9552 8768
rect 9694 8418 9725 8768
rect 9526 8394 9725 8418
rect 14352 8768 14551 8791
rect 14352 8418 14378 8768
rect 14520 8418 14551 8768
rect 14352 8394 14551 8418
rect 19178 8768 19377 8791
rect 19178 8418 19204 8768
rect 19346 8418 19377 8768
rect 19178 8394 19377 8418
rect 24004 8768 24203 8791
rect 24004 8418 24030 8768
rect 24172 8418 24203 8768
rect 24004 8394 24203 8418
rect 18 8372 73 8394
rect 4844 8372 4899 8394
rect 9670 8372 9725 8394
rect 14496 8372 14551 8394
rect 19322 8372 19377 8394
rect 24148 8372 24203 8394
rect 1467 4902 1503 5876
rect 1746 4986 1782 5876
rect 4844 5872 5044 5876
rect 5833 5872 6033 5876
rect 6278 5070 6314 5876
rect 6575 5154 6611 5876
rect 9670 5872 9870 5876
rect 10659 5872 10859 5876
rect 11108 5238 11144 5876
rect 11396 5322 11432 5876
rect 14496 5872 14696 5876
rect 15485 5872 15685 5876
rect 15938 5406 15974 5876
rect 16235 5490 16271 5876
rect 19322 5872 19522 5876
rect 20311 5872 20511 5876
rect 20759 5574 20795 5876
rect 21061 5658 21097 5876
rect 24148 5872 24348 5876
rect 25137 5872 25337 5876
rect 25589 5742 25625 5876
rect 25872 5826 25908 5876
rect 25872 5790 28606 5826
rect 25589 5706 28606 5742
rect 21061 5622 28606 5658
rect 20759 5538 28606 5574
rect 16235 5454 28606 5490
rect 15938 5370 28606 5406
rect 11396 5286 28606 5322
rect 11108 5202 28606 5238
rect 6575 5118 28606 5154
rect 6278 5034 28606 5070
rect 1746 4950 28606 4986
rect 1467 4866 28606 4902
rect 1008 3525 1065 3553
rect 5834 3525 5891 3553
rect 10660 3525 10717 3553
rect 15486 3525 15543 3553
rect 20312 3525 20369 3553
rect 25138 3525 25195 3553
rect 1008 3512 1131 3525
rect 1008 3139 1017 3512
rect 1120 3139 1131 3512
rect 1008 3127 1131 3139
rect 5834 3512 5957 3525
rect 5834 3139 5843 3512
rect 5946 3139 5957 3512
rect 5834 3127 5957 3139
rect 10660 3512 10783 3525
rect 10660 3139 10669 3512
rect 10772 3139 10783 3512
rect 10660 3127 10783 3139
rect 15486 3512 15609 3525
rect 15486 3139 15495 3512
rect 15598 3139 15609 3512
rect 15486 3127 15609 3139
rect 20312 3512 20435 3525
rect 20312 3139 20321 3512
rect 20424 3139 20435 3512
rect 20312 3127 20435 3139
rect 25138 3512 25261 3525
rect 25138 3139 25147 3512
rect 25250 3139 25261 3512
rect 25138 3127 25261 3139
rect 1008 3111 1065 3127
rect 5834 3111 5891 3127
rect 10660 3111 10717 3127
rect 15486 3111 15543 3127
rect 20312 3111 20369 3127
rect 25138 3111 25195 3127
rect 18 2933 24 2952
rect 34 2933 73 2952
rect 18 2925 73 2933
rect 4844 2933 4850 2952
rect 4860 2933 4899 2952
rect 4844 2925 4899 2933
rect 9670 2933 9676 2952
rect 9686 2933 9725 2952
rect 9670 2925 9725 2933
rect 14496 2933 14502 2952
rect 14512 2933 14551 2952
rect 14496 2925 14551 2933
rect 19322 2933 19328 2952
rect 19338 2933 19377 2952
rect 19322 2925 19377 2933
rect 24148 2933 24154 2952
rect 24164 2933 24203 2952
rect 24148 2925 24203 2933
rect -126 2902 73 2925
rect -126 2552 -100 2902
rect 42 2552 73 2902
rect -126 2528 73 2552
rect 4700 2902 4899 2925
rect 4700 2552 4726 2902
rect 4868 2552 4899 2902
rect 4700 2528 4899 2552
rect 9526 2902 9725 2925
rect 9526 2552 9552 2902
rect 9694 2552 9725 2902
rect 9526 2528 9725 2552
rect 14352 2902 14551 2925
rect 14352 2552 14378 2902
rect 14520 2552 14551 2902
rect 14352 2528 14551 2552
rect 19178 2902 19377 2925
rect 19178 2552 19204 2902
rect 19346 2552 19377 2902
rect 19178 2528 19377 2552
rect 24004 2902 24203 2925
rect 24004 2552 24030 2902
rect 24172 2552 24203 2902
rect 24004 2528 24203 2552
rect 18 2506 73 2528
rect 4844 2506 4899 2528
rect 9670 2506 9725 2528
rect 14496 2506 14551 2528
rect 19322 2506 19377 2528
rect 24148 2506 24203 2528
rect 1467 -964 1503 51
rect 1746 -880 1782 75
rect 6278 -796 6314 104
rect 6575 -712 6611 76
rect 11108 -628 11144 72
rect 11396 -544 11432 72
rect 15938 -460 15974 99
rect 16235 -376 16271 49
rect 20759 -292 20795 63
rect 21061 -208 21097 72
rect 25589 -124 25625 72
rect 25872 -40 25908 58
rect 25872 -76 28606 -40
rect 25589 -160 28606 -124
rect 21061 -244 28606 -208
rect 20759 -328 28606 -292
rect 16235 -412 28606 -376
rect 15938 -496 28606 -460
rect 11396 -580 28606 -544
rect 11108 -664 28606 -628
rect 6575 -748 28606 -712
rect 6278 -832 28606 -796
rect 1746 -916 28606 -880
rect 1467 -1000 28606 -964
<< via1 >>
rect 1017 14871 1120 15244
rect 5843 14871 5946 15244
rect 10669 14871 10772 15244
rect 15495 14871 15598 15244
rect 20321 14871 20424 15244
rect 25147 14871 25250 15244
rect -100 14284 42 14634
rect 4726 14284 4868 14634
rect 9552 14284 9694 14634
rect 14378 14284 14520 14634
rect 19204 14284 19346 14634
rect 24030 14284 24172 14634
rect 1017 9005 1120 9378
rect 5843 9005 5946 9378
rect 10669 9005 10772 9378
rect 15495 9005 15598 9378
rect 20321 9005 20424 9378
rect 25147 9005 25250 9378
rect -100 8418 42 8768
rect 4726 8418 4868 8768
rect 9552 8418 9694 8768
rect 14378 8418 14520 8768
rect 19204 8418 19346 8768
rect 24030 8418 24172 8768
rect 1017 3139 1120 3512
rect 5843 3139 5946 3512
rect 10669 3139 10772 3512
rect 15495 3139 15598 3512
rect 20321 3139 20424 3512
rect 25147 3139 25250 3512
rect -100 2552 42 2902
rect 4726 2552 4868 2902
rect 9552 2552 9694 2902
rect 14378 2552 14520 2902
rect 19204 2552 19346 2902
rect 24030 2552 24172 2902
<< metal2 >>
rect 1008 15244 1131 15257
rect 1008 14871 1017 15244
rect 1120 14871 1131 15244
rect 1008 14859 1131 14871
rect -126 14634 64 14657
rect -126 14284 -100 14634
rect 42 14284 64 14634
rect -126 14260 64 14284
rect 1008 9378 1131 9391
rect 1008 9005 1017 9378
rect 1120 9005 1131 9378
rect 1008 8993 1131 9005
rect -126 8768 64 8791
rect -126 8418 -100 8768
rect 42 8418 64 8768
rect -126 8394 64 8418
rect 2661 4630 2861 17164
rect 3693 16362 3893 17200
rect 5834 15244 5957 15257
rect 5834 14871 5843 15244
rect 5946 14871 5957 15244
rect 5834 14859 5957 14871
rect 4700 14634 4890 14657
rect 4700 14284 4726 14634
rect 4868 14284 4890 14634
rect 4700 14260 4890 14284
rect 3693 10183 3893 11318
rect 5834 9378 5957 9391
rect 5834 9005 5843 9378
rect 5946 9005 5957 9378
rect 5834 8993 5957 9005
rect 4700 8768 4890 8791
rect 4700 8418 4726 8768
rect 4868 8418 4890 8768
rect 4700 8394 4890 8418
rect 3693 4317 3893 5483
rect 7487 4317 7687 17164
rect 8519 16362 8719 17188
rect 10660 15244 10783 15257
rect 10660 14871 10669 15244
rect 10772 14871 10783 15244
rect 10660 14859 10783 14871
rect 9526 14634 9716 14657
rect 9526 14284 9552 14634
rect 9694 14284 9716 14634
rect 9526 14260 9716 14284
rect 8519 10183 8719 11306
rect 10660 9378 10783 9391
rect 10660 9005 10669 9378
rect 10772 9005 10783 9378
rect 10660 8993 10783 9005
rect 9526 8768 9716 8791
rect 9526 8418 9552 8768
rect 9694 8418 9716 8768
rect 9526 8394 9716 8418
rect 8519 4317 8719 5459
rect 12313 4317 12513 17164
rect 13345 16362 13545 17212
rect 15486 15244 15609 15257
rect 15486 14871 15495 15244
rect 15598 14871 15609 15244
rect 15486 14859 15609 14871
rect 14352 14634 14542 14657
rect 14352 14284 14378 14634
rect 14520 14284 14542 14634
rect 14352 14260 14542 14284
rect 13345 10183 13545 11330
rect 15486 9378 15609 9391
rect 15486 9005 15495 9378
rect 15598 9005 15609 9378
rect 15486 8993 15609 9005
rect 14352 8768 14542 8791
rect 14352 8418 14378 8768
rect 14520 8418 14542 8768
rect 14352 8394 14542 8418
rect 13345 4317 13545 5459
rect 17139 4317 17339 17164
rect 18171 16049 18371 17212
rect 20312 15244 20435 15257
rect 20312 14871 20321 15244
rect 20424 14871 20435 15244
rect 20312 14859 20435 14871
rect 19178 14634 19368 14657
rect 19178 14284 19204 14634
rect 19346 14284 19368 14634
rect 19178 14260 19368 14284
rect 18171 10183 18371 11330
rect 20312 9378 20435 9391
rect 20312 9005 20321 9378
rect 20424 9005 20435 9378
rect 20312 8993 20435 9005
rect 19178 8768 19368 8791
rect 19178 8418 19204 8768
rect 19346 8418 19368 8768
rect 19178 8394 19368 8418
rect 18171 4317 18371 5459
rect 21965 4317 22165 17164
rect 22997 16049 23197 17188
rect 25138 15244 25261 15257
rect 25138 14871 25147 15244
rect 25250 14871 25261 15244
rect 25138 14859 25261 14871
rect 24004 14634 24194 14657
rect 24004 14284 24030 14634
rect 24172 14284 24194 14634
rect 24004 14260 24194 14284
rect 22997 10183 23197 11318
rect 25138 9378 25261 9391
rect 25138 9005 25147 9378
rect 25250 9005 25261 9378
rect 25138 8993 25261 9005
rect 24004 8768 24194 8791
rect 24004 8418 24030 8768
rect 24172 8418 24194 8768
rect 24004 8394 24194 8418
rect 22997 4317 23197 5483
rect 26791 4317 26991 17164
rect 27823 16049 28023 17200
rect 27823 10183 28023 11330
rect 27823 4317 28023 5447
rect 1008 3512 1131 3525
rect 1008 3139 1017 3512
rect 1120 3139 1131 3512
rect 1008 3127 1131 3139
rect 5834 3512 5957 3525
rect 5834 3139 5843 3512
rect 5946 3139 5957 3512
rect 5834 3127 5957 3139
rect 10660 3512 10783 3525
rect 10660 3139 10669 3512
rect 10772 3139 10783 3512
rect 10660 3127 10783 3139
rect 15486 3512 15609 3525
rect 15486 3139 15495 3512
rect 15598 3139 15609 3512
rect 15486 3127 15609 3139
rect 20312 3512 20435 3525
rect 20312 3139 20321 3512
rect 20424 3139 20435 3512
rect 20312 3127 20435 3139
rect 25138 3512 25261 3525
rect 25138 3139 25147 3512
rect 25250 3139 25261 3512
rect 25138 3127 25261 3139
rect -126 2902 64 2925
rect -126 2552 -100 2902
rect 42 2552 64 2902
rect -126 2528 64 2552
rect 4700 2902 4890 2925
rect 4700 2552 4726 2902
rect 4868 2552 4890 2902
rect 4700 2528 4890 2552
rect 9526 2902 9716 2925
rect 9526 2552 9552 2902
rect 9694 2552 9716 2902
rect 9526 2528 9716 2552
rect 14352 2902 14542 2925
rect 14352 2552 14378 2902
rect 14520 2552 14542 2902
rect 14352 2528 14542 2552
rect 19178 2902 19368 2925
rect 19178 2552 19204 2902
rect 19346 2552 19368 2902
rect 19178 2528 19368 2552
rect 24004 2902 24194 2925
rect 24004 2552 24030 2902
rect 24172 2552 24194 2902
rect 24004 2528 24194 2552
<< via2 >>
rect 1017 14871 1120 15244
rect -100 14284 42 14634
rect 2359 13671 2531 14050
rect 1017 9005 1120 9378
rect -100 8418 42 8768
rect 2359 7805 2531 8184
rect 5843 14871 5946 15244
rect 4726 14284 4868 14634
rect 7185 13671 7357 14050
rect 4024 13069 4202 13449
rect 5843 9005 5946 9378
rect 4726 8418 4868 8768
rect 7185 7805 7357 8184
rect 4024 7203 4202 7583
rect 10669 14871 10772 15244
rect 9552 14284 9694 14634
rect 12011 13671 12183 14050
rect 8850 13069 9028 13449
rect 10669 9005 10772 9378
rect 9552 8418 9694 8768
rect 12011 7805 12183 8184
rect 8850 7203 9028 7583
rect 15495 14871 15598 15244
rect 14378 14284 14520 14634
rect 16837 13671 17009 14050
rect 13676 13069 13854 13449
rect 15495 9005 15598 9378
rect 14378 8418 14520 8768
rect 16837 7805 17009 8184
rect 13676 7203 13854 7583
rect 20321 14871 20424 15244
rect 19204 14284 19346 14634
rect 21663 13671 21835 14050
rect 18502 13069 18680 13449
rect 20321 9005 20424 9378
rect 19204 8418 19346 8768
rect 21663 7805 21835 8184
rect 18502 7203 18680 7583
rect 25147 14871 25250 15244
rect 24030 14284 24172 14634
rect 26489 13671 26661 14050
rect 23328 13069 23506 13449
rect 25147 9005 25250 9378
rect 24030 8418 24172 8768
rect 26489 7805 26661 8184
rect 23328 7203 23506 7583
rect 28154 13069 28332 13449
rect 28154 7203 28332 7583
rect 1017 3139 1120 3512
rect 5843 3139 5946 3512
rect 10669 3139 10772 3512
rect 15495 3139 15598 3512
rect 20321 3139 20424 3512
rect 25147 3139 25250 3512
rect -100 2552 42 2902
rect 4726 2552 4868 2902
rect 9552 2552 9694 2902
rect 14378 2552 14520 2902
rect 19204 2552 19346 2902
rect 24030 2552 24172 2902
rect 2359 1939 2531 2318
rect 7185 1939 7357 2318
rect 12011 1939 12183 2318
rect 16837 1939 17009 2318
rect 21663 1939 21835 2318
rect 26489 1939 26661 2318
rect 4024 1337 4202 1717
rect 8850 1337 9028 1717
rect 13676 1337 13854 1717
rect 18502 1337 18680 1717
rect 23328 1337 23506 1717
rect 28154 1337 28332 1717
<< metal3 >>
rect -77 16971 13561 17171
rect 18127 16971 28595 17171
rect -351 15244 28728 15258
rect -351 14871 1017 15244
rect 1120 14871 5843 15244
rect 5946 15237 10669 15244
rect 10772 15237 15495 15244
rect 5946 14882 10217 15237
rect 10907 14882 15495 15237
rect 5946 14871 10669 14882
rect 10772 14871 15495 14882
rect 15598 14871 20321 15244
rect 20424 14871 25147 15244
rect 25250 14871 28728 15244
rect -351 14858 28728 14871
rect -351 14640 28728 14658
rect -351 14634 15067 14640
rect -351 14284 -100 14634
rect 42 14284 4726 14634
rect 4868 14284 9552 14634
rect 9694 14284 14378 14634
rect 14520 14285 15067 14634
rect 15757 14634 28728 14640
rect 15757 14285 19204 14634
rect 14520 14284 19204 14285
rect 19346 14284 24030 14634
rect 24172 14284 28728 14634
rect -351 14258 28728 14284
rect -351 14050 28728 14058
rect -351 14036 2359 14050
rect -351 13681 581 14036
rect 1271 13681 2359 14036
rect -351 13671 2359 13681
rect 2531 13671 7185 14050
rect 7357 13671 12011 14050
rect 12183 13671 16837 14050
rect 17009 14033 21663 14050
rect 17009 13678 19875 14033
rect 20565 13678 21663 14033
rect 17009 13671 21663 13678
rect 21835 13671 26489 14050
rect 26661 13671 28728 14050
rect -351 13658 28728 13671
rect -351 13449 28728 13458
rect -351 13069 4024 13449
rect 4202 13438 8850 13449
rect 4202 13083 5404 13438
rect 6094 13083 8850 13438
rect 4202 13069 8850 13083
rect 9028 13069 13676 13449
rect 13854 13069 18502 13449
rect 18680 13069 23328 13449
rect 23506 13437 28154 13449
rect 23506 13082 24709 13437
rect 25399 13082 28154 13437
rect 23506 13069 28154 13082
rect 28332 13069 28728 13449
rect -351 13058 28728 13069
rect -76 11105 13562 11305
rect 18126 11105 28594 11305
rect -351 9378 28728 9392
rect -351 9005 1017 9378
rect 1120 9005 5843 9378
rect 5946 9371 10669 9378
rect 10772 9371 15495 9378
rect 5946 9016 10217 9371
rect 10907 9016 15495 9371
rect 5946 9005 10669 9016
rect 10772 9005 15495 9016
rect 15598 9005 20321 9378
rect 20424 9005 25147 9378
rect 25250 9005 28728 9378
rect -351 8992 28728 9005
rect -351 8774 28728 8792
rect -351 8768 15067 8774
rect -351 8418 -100 8768
rect 42 8418 4726 8768
rect 4868 8418 9552 8768
rect 9694 8418 14378 8768
rect 14520 8419 15067 8768
rect 15757 8768 28728 8774
rect 15757 8419 19204 8768
rect 14520 8418 19204 8419
rect 19346 8418 24030 8768
rect 24172 8418 28728 8768
rect -351 8392 28728 8418
rect -351 8184 28728 8192
rect -351 8170 2359 8184
rect -351 7815 581 8170
rect 1271 7815 2359 8170
rect -351 7805 2359 7815
rect 2531 7805 7185 8184
rect 7357 7805 12011 8184
rect 12183 7805 16837 8184
rect 17009 8167 21663 8184
rect 17009 7812 19875 8167
rect 20565 7812 21663 8167
rect 17009 7805 21663 7812
rect 21835 7805 26489 8184
rect 26661 7805 28728 8184
rect -351 7792 28728 7805
rect -351 7583 28728 7592
rect -351 7203 4024 7583
rect 4202 7572 8850 7583
rect 4202 7217 5404 7572
rect 6094 7217 8850 7572
rect 4202 7203 8850 7217
rect 9028 7203 13676 7583
rect 13854 7203 18502 7583
rect 18680 7203 23328 7583
rect 23506 7571 28154 7583
rect 23506 7216 24709 7571
rect 25399 7216 28154 7571
rect 23506 7203 28154 7216
rect 28332 7203 28728 7583
rect -351 7192 28728 7203
rect -77 5239 13561 5439
rect 18127 5239 28595 5439
rect -351 3512 28728 3526
rect -351 3139 1017 3512
rect 1120 3139 5843 3512
rect 5946 3505 10669 3512
rect 10772 3505 15495 3512
rect 5946 3150 10217 3505
rect 10907 3150 15495 3505
rect 5946 3139 10669 3150
rect 10772 3139 15495 3150
rect 15598 3139 20321 3512
rect 20424 3139 25147 3512
rect 25250 3139 28728 3512
rect -351 3126 28728 3139
rect -351 2908 28728 2926
rect -351 2902 15067 2908
rect -351 2552 -100 2902
rect 42 2552 4726 2902
rect 4868 2552 9552 2902
rect 9694 2552 14378 2902
rect 14520 2553 15067 2902
rect 15757 2902 28728 2908
rect 15757 2553 19204 2902
rect 14520 2552 19204 2553
rect 19346 2552 24030 2902
rect 24172 2552 28728 2902
rect -351 2526 28728 2552
rect -351 2318 28728 2326
rect -351 2304 2359 2318
rect -351 1949 581 2304
rect 1271 1949 2359 2304
rect -351 1939 2359 1949
rect 2531 1939 7185 2318
rect 7357 1939 12011 2318
rect 12183 1939 16837 2318
rect 17009 2301 21663 2318
rect 17009 1946 19875 2301
rect 20565 1946 21663 2301
rect 17009 1939 21663 1946
rect 21835 1939 26489 2318
rect 26661 1939 28728 2318
rect -351 1926 28728 1939
rect -351 1717 28728 1726
rect -351 1337 4024 1717
rect 4202 1706 8850 1717
rect 4202 1351 5404 1706
rect 6094 1351 8850 1706
rect 4202 1337 8850 1351
rect 9028 1337 13676 1717
rect 13854 1337 18502 1717
rect 18680 1337 23328 1717
rect 23506 1705 28154 1717
rect 23506 1350 24709 1705
rect 25399 1350 28154 1705
rect 23506 1337 28154 1350
rect 28332 1337 28728 1717
rect -351 1326 28728 1337
<< via3 >>
rect 10217 14882 10669 15237
rect 10669 14882 10772 15237
rect 10772 14882 10907 15237
rect 15067 14285 15757 14640
rect 581 13681 1271 14036
rect 19875 13678 20565 14033
rect 5404 13083 6094 13438
rect 24709 13082 25399 13437
rect 10217 9016 10669 9371
rect 10669 9016 10772 9371
rect 10772 9016 10907 9371
rect 15067 8419 15757 8774
rect 581 7815 1271 8170
rect 19875 7812 20565 8167
rect 5404 7217 6094 7572
rect 24709 7216 25399 7571
rect 10217 3150 10669 3505
rect 10669 3150 10772 3505
rect 10772 3150 10907 3505
rect 15067 2553 15757 2908
rect 581 1949 1271 2304
rect 19875 1946 20565 2301
rect 5404 1351 6094 1706
rect 24709 1350 25399 1705
<< metal4 >>
rect 558 14036 1297 17274
rect 558 13681 581 14036
rect 1271 13681 1297 14036
rect 558 8170 1297 13681
rect 558 7815 581 8170
rect 1271 7815 1297 8170
rect 558 2304 1297 7815
rect 558 1949 581 2304
rect 1271 1949 1297 2304
rect 558 -599 1297 1949
rect 5384 13438 6123 17274
rect 5384 13083 5404 13438
rect 6094 13083 6123 13438
rect 5384 7572 6123 13083
rect 5384 7217 5404 7572
rect 6094 7217 6123 7572
rect 5384 1706 6123 7217
rect 5384 1351 5404 1706
rect 6094 1351 6123 1706
rect 5384 -599 6123 1351
rect 10210 15237 10949 17274
rect 10210 14882 10217 15237
rect 10907 14882 10949 15237
rect 10210 9371 10949 14882
rect 10210 9016 10217 9371
rect 10907 9016 10949 9371
rect 10210 3505 10949 9016
rect 10210 3150 10217 3505
rect 10907 3150 10949 3505
rect 10210 -599 10949 3150
rect 15036 14640 15775 17274
rect 15036 14285 15067 14640
rect 15757 14285 15775 14640
rect 15036 8774 15775 14285
rect 15036 8419 15067 8774
rect 15757 8419 15775 8774
rect 15036 2908 15775 8419
rect 15036 2553 15067 2908
rect 15757 2553 15775 2908
rect 15036 -599 15775 2553
rect 19862 14033 20601 17274
rect 19862 13678 19875 14033
rect 20565 13678 20601 14033
rect 19862 8167 20601 13678
rect 19862 7812 19875 8167
rect 20565 7812 20601 8167
rect 19862 2301 20601 7812
rect 19862 1946 19875 2301
rect 20565 1946 20601 2301
rect 19862 -599 20601 1946
rect 24688 13437 25427 17274
rect 24688 13082 24709 13437
rect 25399 13082 25427 13437
rect 24688 7571 25427 13082
rect 24688 7216 24709 7571
rect 25399 7216 25427 7571
rect 24688 1705 25427 7216
rect 24688 1350 24709 1705
rect 25399 1350 25427 1705
rect 24688 -599 25427 1350
use cv3_via2_36cut  cv3_via2_36cut_0
timestamp 1719173892
transform 1 0 -542238 0 1 -86992
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_1
timestamp 1719173892
transform 1 0 -527772 0 1 -87028
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_2
timestamp 1719173892
transform 1 0 -547012 0 1 -87020
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_3
timestamp 1719173892
transform 1 0 -551878 0 1 -87001
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_4
timestamp 1719173892
transform 1 0 -537355 0 1 -87010
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_5
timestamp 1719173892
transform 1 0 -532573 0 1 -87028
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_6
timestamp 1719173892
transform 1 0 -527772 0 1 -75296
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_7
timestamp 1719173892
transform 1 0 -532573 0 1 -75296
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_8
timestamp 1719173892
transform 1 0 -537355 0 1 -75278
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_9
timestamp 1719173892
transform 1 0 -551878 0 1 -75269
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_10
timestamp 1719173892
transform 1 0 -542238 0 1 -75260
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_11
timestamp 1719173892
transform 1 0 -547012 0 1 -75288
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_12
timestamp 1719173892
transform 1 0 -551878 0 1 -81135
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_13
timestamp 1719173892
transform 1 0 -547012 0 1 -81154
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_14
timestamp 1719173892
transform 1 0 -542238 0 1 -81126
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_15
timestamp 1719173892
transform 1 0 -537355 0 1 -81144
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_16
timestamp 1719173892
transform 1 0 -532573 0 1 -81162
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_17
timestamp 1719173892
transform 1 0 -527772 0 1 -81162
box 555256 92202 556228 92502
use isolated_switch_large  isolated_switch_large_0 ../dependencies/sky130_ef_ip__analog_switches/mag
array 0 2 5866 0 5 -4826
timestamp 1719093964
transform 0 -1 1336 1 0 -656
box 660 -3110 5486 1338
<< labels >>
flabel metal2 2661 16964 2861 17164 0 FreeSans 1120 0 0 0 ulpcomp_n
flabel metal2 7487 16964 7687 17164 0 FreeSans 1120 0 0 0 comp_n
flabel metal2 12313 16964 12513 17164 0 FreeSans 1120 0 0 0 adc1
flabel metal2 17139 16964 17339 17164 0 FreeSans 1120 0 0 0 ulpcomp_p
flabel metal2 21965 16964 22165 17164 0 FreeSans 1120 0 0 0 comp_p
flabel metal2 26791 16964 26991 17164 0 FreeSans 1120 0 0 0 adc0
flabel metal3 28435 11105 28594 11205 0 FreeSans 1120 0 0 0 left_hgbw_opamp_out
flabel metal3 28380 16971 28595 17171 0 FreeSans 1120 0 0 0 left_instramp_out
flabel metal3 -76 5239 124 5439 0 FreeSans 1120 0 0 0 left_lp_opamp_out
flabel metal3 -76 11105 124 11305 0 FreeSans 1120 0 0 0 right_hgbw_opamp_out
flabel metal3 -76 16971 124 17171 0 FreeSans 1120 0 0 0 right_instramp_out
flabel metal3 28395 5239 28595 5439 0 FreeSans 1120 0 0 0 right_lp_opamp_out
flabel metal4 894 -346 894 -346 0 FreeSans 1280 0 0 0 avdd
flabel metal4 5718 -362 5718 -362 0 FreeSans 1280 0 0 0 avss
flabel metal4 10558 -362 10558 -362 0 FreeSans 1280 0 0 0 dvdd
flabel metal4 15376 -342 15376 -342 0 FreeSans 1280 0 0 0 dvss
<< end >>
