magic
tech sky130A
magscale 1 2
timestamp 1724447141
<< metal1 >>
rect 12895 19350 12901 19357
rect -648 19314 12901 19350
rect 12895 19305 12901 19314
rect 12953 19305 12959 19357
rect 17423 19306 17429 19358
rect 17481 19350 17487 19358
rect 17481 19314 26691 19350
rect 17481 19306 17487 19314
rect 8408 19266 8414 19272
rect -648 19230 8414 19266
rect 8408 19220 8414 19230
rect 8466 19220 8472 19272
rect 21950 19222 21956 19274
rect 22008 19266 22014 19274
rect 22008 19230 26691 19266
rect 22008 19222 22014 19230
rect 3871 19182 3877 19185
rect -648 19146 3877 19182
rect 3871 19133 3877 19146
rect 3929 19133 3935 19185
rect 26462 19138 26468 19190
rect 26520 19182 26526 19190
rect 26520 19146 26691 19182
rect 26520 19138 26526 19146
rect 2782 19021 3474 19038
rect 2782 19008 2809 19021
rect 2781 18860 2809 19008
rect 2782 18838 2809 18860
rect 3440 18838 3474 19021
rect 7298 19021 7990 19038
rect 7298 19008 7325 19021
rect 7297 18860 7325 19008
rect 2782 18822 3474 18838
rect 7298 18838 7325 18860
rect 7956 18838 7990 19021
rect 11814 19021 12506 19038
rect 11814 19008 11841 19021
rect 11813 18860 11841 19008
rect 7298 18822 7990 18838
rect 11814 18838 11841 18860
rect 12472 18838 12506 19021
rect 16330 19021 17022 19038
rect 16330 19008 16357 19021
rect 16329 18860 16357 19008
rect 11814 18822 12506 18838
rect 16330 18838 16357 18860
rect 16988 18838 17022 19021
rect 20846 19021 21538 19038
rect 20846 19008 20873 19021
rect 20845 18860 20873 19008
rect 16330 18822 17022 18838
rect 20846 18838 20873 18860
rect 21504 18838 21538 19021
rect 25362 19021 26054 19038
rect 25362 19008 25389 19021
rect 25361 18860 25389 19008
rect 20846 18822 21538 18838
rect 25362 18838 25389 18860
rect 26020 18838 26054 19021
rect 25362 18822 26054 18838
rect 3243 18215 3651 18251
rect 3243 17945 3278 18215
rect 3614 17945 3651 18215
rect 3243 17908 3651 17945
rect 7759 18215 8167 18251
rect 7759 17945 7794 18215
rect 8130 17945 8167 18215
rect 7759 17908 8167 17945
rect 12275 18215 12683 18251
rect 12275 17945 12310 18215
rect 12646 17945 12683 18215
rect 12275 17908 12683 17945
rect 16791 18215 17199 18251
rect 16791 17945 16826 18215
rect 17162 17945 17199 18215
rect 16791 17908 17199 17945
rect 21307 18215 21715 18251
rect 21307 17945 21342 18215
rect 21678 17945 21715 18215
rect 21307 17908 21715 17945
rect 25823 18215 26231 18251
rect 25823 17945 25858 18215
rect 26194 17945 26231 18215
rect 25823 17908 26231 17945
rect 3871 17487 3877 17496
rect 3422 17451 3877 17487
rect 3871 17444 3877 17451
rect 3929 17444 3935 17496
rect 8408 17485 8414 17491
rect 7945 17449 8414 17485
rect 8408 17439 8414 17449
rect 8466 17439 8472 17491
rect 12895 17484 12901 17492
rect 12488 17448 12901 17484
rect 12895 17440 12901 17448
rect 12953 17440 12959 17492
rect 26462 17485 26468 17493
rect 17423 17477 17429 17485
rect 16985 17441 17429 17477
rect 17423 17433 17429 17441
rect 17481 17433 17487 17485
rect 21950 17476 21956 17484
rect 21481 17440 21956 17476
rect 21950 17432 21956 17440
rect 22008 17432 22014 17484
rect 26029 17449 26468 17485
rect 26462 17441 26468 17449
rect 26520 17441 26526 17493
rect 12903 14717 12909 14725
rect -648 14681 12909 14717
rect 12903 14673 12909 14681
rect 12961 14673 12967 14725
rect 17401 14673 17407 14725
rect 17459 14717 17465 14725
rect 17459 14681 26780 14717
rect 17459 14673 17465 14681
rect 8402 14633 8408 14641
rect -648 14597 8408 14633
rect 8402 14589 8408 14597
rect 8460 14589 8466 14641
rect 21945 14589 21951 14641
rect 22003 14633 22009 14641
rect 22003 14597 26780 14633
rect 22003 14589 22009 14597
rect 3871 14549 3877 14557
rect -648 14513 3877 14549
rect 3871 14505 3877 14513
rect 3929 14505 3935 14557
rect 26489 14505 26495 14557
rect 26547 14549 26553 14557
rect 26547 14513 26780 14549
rect 26547 14505 26553 14513
rect 2782 14388 3474 14405
rect 2782 14375 2809 14388
rect 2781 14227 2809 14375
rect 2782 14205 2809 14227
rect 3440 14205 3474 14388
rect 7298 14388 7990 14405
rect 7298 14375 7325 14388
rect 7297 14227 7325 14375
rect 2782 14189 3474 14205
rect 7298 14205 7325 14227
rect 7956 14205 7990 14388
rect 11814 14388 12506 14405
rect 11814 14375 11841 14388
rect 11813 14227 11841 14375
rect 7298 14189 7990 14205
rect 11814 14205 11841 14227
rect 12472 14205 12506 14388
rect 16330 14388 17022 14405
rect 16330 14375 16357 14388
rect 16329 14227 16357 14375
rect 11814 14189 12506 14205
rect 16330 14205 16357 14227
rect 16988 14205 17022 14388
rect 20846 14388 21538 14405
rect 20846 14375 20873 14388
rect 20845 14227 20873 14375
rect 16330 14189 17022 14205
rect 20846 14205 20873 14227
rect 21504 14205 21538 14388
rect 25362 14388 26054 14405
rect 25362 14375 25389 14388
rect 25361 14227 25389 14375
rect 20846 14189 21538 14205
rect 25362 14205 25389 14227
rect 26020 14205 26054 14388
rect 25362 14189 26054 14205
rect 3243 13582 3651 13618
rect 3243 13312 3278 13582
rect 3614 13312 3651 13582
rect 3243 13275 3651 13312
rect 7759 13582 8167 13618
rect 7759 13312 7794 13582
rect 8130 13312 8167 13582
rect 7759 13275 8167 13312
rect 12275 13582 12683 13618
rect 12275 13312 12310 13582
rect 12646 13312 12683 13582
rect 12275 13275 12683 13312
rect 16791 13582 17199 13618
rect 16791 13312 16826 13582
rect 17162 13312 17199 13582
rect 16791 13275 17199 13312
rect 21307 13582 21715 13618
rect 21307 13312 21342 13582
rect 21678 13312 21715 13582
rect 21307 13275 21715 13312
rect 25823 13582 26231 13618
rect 25823 13312 25858 13582
rect 26194 13312 26231 13582
rect 25823 13275 26231 13312
rect 12903 12856 12909 12862
rect 3871 12847 3877 12855
rect 3423 12811 3877 12847
rect 3871 12803 3877 12811
rect 3929 12803 3935 12855
rect 8402 12841 8408 12849
rect 7939 12805 8408 12841
rect 8402 12797 8408 12805
rect 8460 12797 8466 12849
rect 12476 12820 12909 12856
rect 12903 12810 12909 12820
rect 12961 12810 12967 12862
rect 17401 12848 17407 12856
rect 16952 12812 17407 12848
rect 17401 12804 17407 12812
rect 17459 12804 17465 12856
rect 21945 12849 21951 12857
rect 21476 12813 21951 12849
rect 21945 12805 21951 12813
rect 22003 12805 22009 12857
rect 26489 12848 26495 12856
rect 26020 12812 26495 12848
rect 26489 12804 26495 12812
rect 26547 12804 26553 12856
rect 26172 10221 26959 10257
rect 12914 10084 12920 10092
rect -648 10048 12920 10084
rect 12914 10040 12920 10048
rect 12972 10040 12978 10092
rect 17426 10040 17432 10092
rect 17484 10084 17490 10092
rect 26172 10084 26208 10221
rect 17484 10048 26208 10084
rect 26256 10137 26959 10173
rect 17484 10040 17490 10048
rect 8396 10000 8402 10008
rect -648 9964 8402 10000
rect 8396 9956 8402 9964
rect 8454 9956 8460 10008
rect 21938 9956 21944 10008
rect 21996 10000 22002 10008
rect 26256 10000 26292 10137
rect 26403 10045 26409 10097
rect 26461 10089 26467 10097
rect 26461 10053 26959 10089
rect 26461 10045 26467 10053
rect 21996 9964 26292 10000
rect 21996 9956 22002 9964
rect 3863 9916 3869 9924
rect -648 9880 3869 9916
rect 3863 9872 3869 9880
rect 3921 9872 3927 9924
rect 26501 9887 26507 9939
rect 26559 9931 26565 9939
rect 26559 9895 26959 9931
rect 26559 9887 26565 9895
rect 2782 9755 3474 9772
rect 2782 9572 2809 9755
rect 3440 9572 3474 9755
rect 7298 9755 7990 9772
rect 7298 9742 7325 9755
rect 7297 9594 7325 9742
rect 2782 9556 3474 9572
rect 7298 9572 7325 9594
rect 7956 9572 7990 9755
rect 11814 9755 12506 9772
rect 11814 9742 11841 9755
rect 11813 9594 11841 9742
rect 7298 9556 7990 9572
rect 11814 9572 11841 9594
rect 12472 9572 12506 9755
rect 16330 9755 17022 9772
rect 16330 9742 16357 9755
rect 16329 9594 16357 9742
rect 11814 9556 12506 9572
rect 16330 9572 16357 9594
rect 16988 9572 17022 9755
rect 20846 9755 21538 9772
rect 20846 9742 20873 9755
rect 20845 9594 20873 9742
rect 16330 9556 17022 9572
rect 20846 9572 20873 9594
rect 21504 9572 21538 9755
rect 25362 9755 26054 9772
rect 25362 9742 25389 9755
rect 25361 9594 25389 9742
rect 20846 9556 21538 9572
rect 25362 9572 25389 9594
rect 26020 9572 26054 9755
rect 29878 9755 30570 9772
rect 29878 9742 29905 9755
rect 29877 9594 29905 9742
rect 25362 9556 26054 9572
rect 29878 9572 29905 9594
rect 30536 9572 30570 9755
rect 34394 9755 35086 9772
rect 34394 9742 34421 9755
rect 34393 9594 34421 9742
rect 29878 9556 30570 9572
rect 34394 9572 34421 9594
rect 35052 9572 35086 9755
rect 38910 9755 39602 9772
rect 38910 9742 38937 9755
rect 38909 9594 38937 9742
rect 34394 9556 35086 9572
rect 38910 9572 38937 9594
rect 39568 9572 39602 9755
rect 43426 9755 44118 9772
rect 43426 9742 43453 9755
rect 43425 9594 43453 9742
rect 38910 9556 39602 9572
rect 43426 9572 43453 9594
rect 44084 9572 44118 9755
rect 43426 9556 44118 9572
rect 3243 9089 3511 9125
rect 3243 8679 3278 9089
rect 3474 8679 3511 9089
rect 3243 8642 3511 8679
rect 7759 9089 8027 9125
rect 7759 8679 7794 9089
rect 7990 8679 8027 9089
rect 7759 8642 8027 8679
rect 12275 9089 12543 9124
rect 12275 8679 12310 9089
rect 12506 8679 12543 9089
rect 12275 8642 12543 8679
rect 16791 9089 17059 9125
rect 16791 8679 16826 9089
rect 17022 8679 17059 9089
rect 16791 8642 17059 8679
rect 21307 9089 21575 9125
rect 21307 8679 21342 9089
rect 21538 8679 21575 9089
rect 21307 8642 21575 8679
rect 25823 9089 26091 9125
rect 25823 8679 25858 9089
rect 26054 8679 26091 9089
rect 39371 9089 39639 9125
rect 25823 8642 26091 8679
rect 30339 8949 30747 8985
rect 30339 8679 30374 8949
rect 30710 8679 30747 8949
rect 30339 8642 30747 8679
rect 34855 8949 35263 8985
rect 34855 8679 34890 8949
rect 35226 8679 35263 8949
rect 34855 8642 35263 8679
rect 39371 8679 39406 9089
rect 39602 8679 39639 9089
rect 39371 8642 39639 8679
rect 43887 9089 44155 9125
rect 43887 8679 43922 9089
rect 44118 8679 44155 9089
rect 43887 8642 44155 8679
rect 35435 8229 35441 8237
rect 3863 8216 3869 8224
rect 3428 8180 3869 8216
rect 3863 8172 3869 8180
rect 3921 8172 3927 8224
rect 8396 8210 8402 8218
rect 7959 8174 8402 8210
rect 8396 8166 8402 8174
rect 8454 8166 8460 8218
rect 12914 8216 12920 8224
rect 12442 8180 12920 8216
rect 12914 8172 12920 8180
rect 12972 8172 12978 8224
rect 17426 8219 17432 8227
rect 16971 8183 17432 8219
rect 17426 8175 17432 8183
rect 17484 8175 17490 8227
rect 21938 8219 21944 8227
rect 21493 8183 21944 8219
rect 21938 8175 21944 8183
rect 21996 8175 22002 8227
rect 26403 8216 26409 8224
rect 25999 8180 26409 8216
rect 26403 8172 26409 8180
rect 26461 8172 26467 8224
rect 30924 8216 30930 8224
rect 30555 8180 30930 8216
rect 30924 8172 30930 8180
rect 30982 8172 30988 8224
rect 35040 8193 35441 8229
rect 35435 8185 35441 8193
rect 35493 8185 35499 8237
rect 39662 8221 39669 8233
rect 39581 8193 39669 8221
rect 39662 8181 39669 8193
rect 39721 8221 39727 8233
rect 39721 8193 39733 8221
rect 39721 8181 39727 8193
rect 40382 7883 40388 7935
rect 40440 7923 40446 7935
rect 44072 7923 44100 8214
rect 40440 7895 44100 7923
rect 40440 7883 40446 7895
rect 12894 5451 12900 5459
rect -648 5415 12900 5451
rect 12894 5407 12900 5415
rect 12952 5407 12958 5459
rect 17439 5407 17445 5459
rect 17497 5451 17503 5459
rect 26501 5451 26507 5459
rect 17497 5415 26507 5451
rect 17497 5407 17503 5415
rect 26501 5407 26507 5415
rect 26559 5407 26565 5459
rect 31017 5375 31069 5381
rect 8397 5367 8403 5375
rect -648 5331 8403 5367
rect 8397 5323 8403 5331
rect 8455 5323 8461 5375
rect 21952 5323 21958 5375
rect 22010 5367 22016 5375
rect 22010 5331 31017 5367
rect 22010 5323 22016 5331
rect 31017 5317 31069 5323
rect 3864 5283 3870 5291
rect -648 5247 3870 5283
rect 3864 5239 3870 5247
rect 3922 5239 3928 5291
rect 26415 5239 26421 5291
rect 26473 5283 26479 5291
rect 35539 5283 35545 5291
rect 26473 5247 35545 5283
rect 26473 5239 26479 5247
rect 35539 5239 35545 5247
rect 35597 5239 35603 5291
rect 2782 5122 3474 5139
rect 2782 5109 2809 5122
rect 2781 4961 2809 5109
rect 2782 4939 2809 4961
rect 3440 4939 3474 5122
rect 7298 5122 7990 5139
rect 7298 5109 7325 5122
rect 7297 4961 7325 5109
rect 2782 4923 3474 4939
rect 7298 4939 7325 4961
rect 7956 4939 7990 5122
rect 11814 5122 12506 5139
rect 11814 5109 11841 5122
rect 11813 4961 11841 5109
rect 7298 4923 7990 4939
rect 11814 4939 11841 4961
rect 12472 4939 12506 5122
rect 16330 5122 17022 5139
rect 16330 5109 16357 5122
rect 16329 4961 16357 5109
rect 11814 4923 12506 4939
rect 16330 4939 16357 4961
rect 16988 4939 17022 5122
rect 20846 5122 21538 5139
rect 20846 5109 20873 5122
rect 20845 4961 20873 5109
rect 16330 4923 17022 4939
rect 20846 4939 20873 4961
rect 21504 4939 21538 5122
rect 25362 5122 26054 5139
rect 25362 5109 25389 5122
rect 25361 4961 25389 5109
rect 20846 4923 21538 4939
rect 25362 4939 25389 4961
rect 26020 4939 26054 5122
rect 29878 5122 30570 5139
rect 29878 5109 29905 5122
rect 29877 4961 29905 5109
rect 25362 4923 26054 4939
rect 29878 4939 29905 4961
rect 30536 4939 30570 5122
rect 34394 5122 35086 5139
rect 34394 5109 34421 5122
rect 34393 4961 34421 5109
rect 29878 4923 30570 4939
rect 34394 4939 34421 4961
rect 35052 4939 35086 5122
rect 38910 5122 39602 5139
rect 38910 5109 38937 5122
rect 38909 4961 38937 5109
rect 34394 4923 35086 4939
rect 38910 4939 38937 4961
rect 39568 4939 39602 5122
rect 43426 5122 44118 5139
rect 43426 5109 43453 5122
rect 43425 4961 43453 5109
rect 38910 4923 39602 4939
rect 43426 4939 43453 4961
rect 44084 4939 44118 5122
rect 43426 4923 44118 4939
rect 3243 4456 3511 4492
rect 3243 4046 3278 4456
rect 3474 4046 3511 4456
rect 3243 4009 3511 4046
rect 7759 4456 8027 4492
rect 7759 4046 7794 4456
rect 7990 4046 8027 4456
rect 7759 4009 8027 4046
rect 12275 4456 12543 4492
rect 12275 4046 12310 4456
rect 12506 4046 12543 4456
rect 12275 4009 12543 4046
rect 16791 4456 17059 4491
rect 16791 4046 16826 4456
rect 17022 4046 17059 4456
rect 16791 4009 17059 4046
rect 21307 4456 21575 4492
rect 21307 4046 21342 4456
rect 21538 4046 21575 4456
rect 21307 4009 21575 4046
rect 25823 4456 26091 4492
rect 25823 4046 25858 4456
rect 26054 4046 26091 4456
rect 43887 4456 44155 4492
rect 25823 4009 26091 4046
rect 30339 4316 30747 4352
rect 30339 4046 30374 4316
rect 30710 4046 30747 4316
rect 30339 4009 30747 4046
rect 34855 4316 35263 4352
rect 34855 4046 34890 4316
rect 35226 4046 35263 4316
rect 34855 4009 35263 4046
rect 39371 4316 39779 4352
rect 39371 4046 39406 4316
rect 39742 4046 39779 4316
rect 39371 4009 39779 4046
rect 43887 4046 43922 4456
rect 44118 4046 44155 4456
rect 43887 4009 44155 4046
rect 8397 3585 8403 3593
rect 3864 3576 3870 3584
rect 3439 3540 3870 3576
rect 3864 3532 3870 3540
rect 3922 3532 3928 3584
rect 7962 3549 8403 3585
rect 8397 3541 8403 3549
rect 8455 3541 8461 3593
rect 12894 3585 12900 3593
rect 12462 3549 12900 3585
rect 12894 3541 12900 3549
rect 12952 3541 12958 3593
rect 26415 3587 26421 3595
rect 17439 3577 17445 3585
rect 16983 3541 17445 3577
rect 17439 3533 17445 3541
rect 17497 3533 17503 3585
rect 21952 3577 21958 3585
rect 21499 3541 21958 3577
rect 21952 3533 21958 3541
rect 22010 3533 22016 3585
rect 26037 3551 26421 3587
rect 26415 3543 26421 3551
rect 26473 3543 26479 3595
rect 39967 3580 39973 3592
rect 30516 3537 30669 3573
rect 30633 837 30669 3537
rect 35040 3529 35167 3565
rect 39532 3552 39973 3580
rect 39967 3540 39973 3552
rect 40025 3540 40031 3592
rect -599 801 30671 837
rect 30924 753 30930 764
rect -599 717 30930 753
rect 30924 712 30930 717
rect 30982 712 30988 764
rect 35131 669 35167 3529
rect 40045 3251 40051 3303
rect 40103 3291 40109 3303
rect 44084 3291 44112 3613
rect 40103 3263 44112 3291
rect 40103 3251 40109 3263
rect -599 633 35167 669
rect 35435 585 35441 591
rect -599 549 35441 585
rect 35435 539 35441 549
rect 35493 539 35499 591
<< via1 >>
rect 12901 19305 12953 19357
rect 17429 19306 17481 19358
rect 8414 19220 8466 19272
rect 21956 19222 22008 19274
rect 3877 19133 3929 19185
rect 26468 19138 26520 19190
rect 2809 18838 3440 19021
rect 7325 18838 7956 19021
rect 11841 18838 12472 19021
rect 16357 18838 16988 19021
rect 20873 18838 21504 19021
rect 25389 18838 26020 19021
rect 3278 17945 3614 18215
rect 7794 17945 8130 18215
rect 12310 17945 12646 18215
rect 16826 17945 17162 18215
rect 21342 17945 21678 18215
rect 25858 17945 26194 18215
rect 3877 17444 3929 17496
rect 8414 17439 8466 17491
rect 12901 17440 12953 17492
rect 17429 17433 17481 17485
rect 21956 17432 22008 17484
rect 26468 17441 26520 17493
rect 12909 14673 12961 14725
rect 17407 14673 17459 14725
rect 8408 14589 8460 14641
rect 21951 14589 22003 14641
rect 3877 14505 3929 14557
rect 26495 14505 26547 14557
rect 2809 14205 3440 14388
rect 7325 14205 7956 14388
rect 11841 14205 12472 14388
rect 16357 14205 16988 14388
rect 20873 14205 21504 14388
rect 25389 14205 26020 14388
rect 3278 13312 3614 13582
rect 7794 13312 8130 13582
rect 12310 13312 12646 13582
rect 16826 13312 17162 13582
rect 21342 13312 21678 13582
rect 25858 13312 26194 13582
rect 3877 12803 3929 12855
rect 8408 12797 8460 12849
rect 12909 12810 12961 12862
rect 17407 12804 17459 12856
rect 21951 12805 22003 12857
rect 26495 12804 26547 12856
rect 12920 10040 12972 10092
rect 17432 10040 17484 10092
rect 8402 9956 8454 10008
rect 21944 9956 21996 10008
rect 26409 10045 26461 10097
rect 3869 9872 3921 9924
rect 26507 9887 26559 9939
rect 2809 9572 3440 9755
rect 7325 9572 7956 9755
rect 11841 9572 12472 9755
rect 16357 9572 16988 9755
rect 20873 9572 21504 9755
rect 25389 9572 26020 9755
rect 29905 9572 30536 9755
rect 34421 9572 35052 9755
rect 38937 9572 39568 9755
rect 43453 9572 44084 9755
rect 3278 8679 3474 9089
rect 7794 8679 7990 9089
rect 12310 8679 12506 9089
rect 16826 8679 17022 9089
rect 21342 8679 21538 9089
rect 25858 8679 26054 9089
rect 30374 8679 30710 8949
rect 34890 8679 35226 8949
rect 39406 8679 39602 9089
rect 43922 8679 44118 9089
rect 3869 8172 3921 8224
rect 8402 8166 8454 8218
rect 12920 8172 12972 8224
rect 17432 8175 17484 8227
rect 21944 8175 21996 8227
rect 26409 8172 26461 8224
rect 30930 8172 30982 8224
rect 35441 8185 35493 8237
rect 39669 8181 39721 8233
rect 40388 7883 40440 7935
rect 12900 5407 12952 5459
rect 17445 5407 17497 5459
rect 26507 5407 26559 5459
rect 8403 5323 8455 5375
rect 21958 5323 22010 5375
rect 31017 5323 31069 5375
rect 3870 5239 3922 5291
rect 26421 5239 26473 5291
rect 35545 5239 35597 5291
rect 2809 4939 3440 5122
rect 7325 4939 7956 5122
rect 11841 4939 12472 5122
rect 16357 4939 16988 5122
rect 20873 4939 21504 5122
rect 25389 4939 26020 5122
rect 29905 4939 30536 5122
rect 34421 4939 35052 5122
rect 38937 4939 39568 5122
rect 43453 4939 44084 5122
rect 3278 4046 3474 4456
rect 7794 4046 7990 4456
rect 12310 4046 12506 4456
rect 16826 4046 17022 4456
rect 21342 4046 21538 4456
rect 25858 4046 26054 4456
rect 30374 4046 30710 4316
rect 34890 4046 35226 4316
rect 39406 4046 39742 4316
rect 43922 4046 44118 4456
rect 3870 3532 3922 3584
rect 8403 3541 8455 3593
rect 12900 3541 12952 3593
rect 17445 3533 17497 3585
rect 21958 3533 22010 3585
rect 26421 3543 26473 3595
rect 39973 3540 40025 3592
rect 30930 712 30982 764
rect 40051 3251 40103 3303
rect 35441 539 35493 591
<< metal2 >>
rect 12901 19357 12953 19363
rect 12901 19299 12953 19305
rect 17429 19358 17481 19364
rect 17429 19300 17481 19306
rect 8414 19272 8466 19278
rect 8414 19214 8466 19220
rect 3877 19185 3929 19191
rect 3877 19127 3929 19133
rect 2781 19021 3473 19038
rect 2781 18838 2809 19021
rect 3440 18838 3473 19021
rect 2781 18822 3473 18838
rect 3243 18215 3651 18251
rect 3243 17945 3278 18215
rect 3614 17945 3651 18215
rect 3243 17908 3651 17945
rect 3885 17502 3921 19127
rect 7297 19021 7989 19038
rect 7297 18838 7325 19021
rect 7956 18838 7989 19021
rect 7297 18822 7989 18838
rect 7759 18215 8167 18251
rect 7759 17945 7794 18215
rect 8130 17945 8167 18215
rect 7759 17908 8167 17945
rect 3877 17496 3929 17502
rect 8422 17497 8458 19214
rect 11813 19021 12505 19038
rect 11813 18838 11841 19021
rect 12472 18838 12505 19021
rect 11813 18822 12505 18838
rect 12275 18215 12683 18251
rect 12275 17945 12310 18215
rect 12646 17945 12683 18215
rect 12275 17908 12683 17945
rect 12909 17498 12945 19299
rect 16329 19021 17021 19038
rect 16329 18838 16357 19021
rect 16988 18838 17021 19021
rect 16329 18822 17021 18838
rect 16791 18215 17199 18251
rect 16791 17945 16826 18215
rect 17162 17945 17199 18215
rect 16791 17908 17199 17945
rect 3877 17438 3929 17444
rect 8414 17491 8466 17497
rect 8414 17433 8466 17439
rect 12901 17492 12953 17498
rect 17437 17491 17473 19300
rect 21956 19274 22008 19280
rect 21956 19216 22008 19222
rect 20845 19021 21537 19038
rect 20845 18838 20873 19021
rect 21504 18838 21537 19021
rect 20845 18822 21537 18838
rect 21307 18215 21715 18251
rect 21307 17945 21342 18215
rect 21678 17945 21715 18215
rect 21307 17908 21715 17945
rect 12901 17434 12953 17440
rect 17429 17485 17481 17491
rect 21964 17490 22000 19216
rect 26468 19190 26520 19196
rect 26468 19132 26520 19138
rect 25361 19021 26053 19038
rect 25361 18838 25389 19021
rect 26020 18838 26053 19021
rect 25361 18822 26053 18838
rect 25823 18215 26231 18251
rect 25823 17945 25858 18215
rect 26194 17945 26231 18215
rect 25823 17908 26231 17945
rect 26476 17499 26512 19132
rect 26468 17493 26520 17499
rect 17429 17427 17481 17433
rect 21956 17484 22008 17490
rect 26468 17435 26520 17441
rect 21956 17426 22008 17432
rect 4030 16352 4166 16386
rect 8546 16352 8682 16362
rect 13062 16352 13198 16370
rect 17578 16352 17714 16362
rect 22094 16352 22230 16378
rect -318 16346 50 16352
rect -492 15920 50 16346
rect 4030 15920 4548 16352
rect 8546 15920 9024 16352
rect 13062 15920 13542 16352
rect 17578 15920 18052 16352
rect 22094 15920 22586 16352
rect -492 7086 -356 15920
rect 3877 14557 3929 14563
rect 3877 14499 3929 14505
rect 2781 14388 3473 14405
rect 2781 14205 2809 14388
rect 3440 14205 3473 14388
rect 2781 14189 3473 14205
rect 3243 13582 3651 13618
rect 3243 13312 3278 13582
rect 3614 13312 3651 13582
rect 3243 13275 3651 13312
rect 3885 12861 3921 14499
rect 3877 12855 3929 12861
rect 3877 12797 3929 12803
rect 3630 11719 3766 11759
rect 3030 11287 3766 11719
rect 2781 9755 3473 9772
rect 2781 9572 2809 9755
rect 3440 9572 3473 9755
rect 2781 9555 3473 9572
rect 3243 9089 3511 9125
rect 3243 8679 3278 9089
rect 3474 8679 3511 9089
rect 3243 8642 3511 8679
rect -492 6654 34 7086
rect -492 1342 -356 6654
rect 2781 5122 3473 5139
rect 2781 4939 2809 5122
rect 3440 4939 3473 5122
rect 2781 4923 3473 4939
rect 3243 4456 3511 4492
rect 3243 4046 3278 4456
rect 3474 4046 3511 4456
rect 3243 4009 3511 4046
rect 3630 2453 3766 11287
rect 3869 9924 3921 9930
rect 3869 9866 3921 9872
rect 3877 8230 3913 9866
rect 3869 8224 3921 8230
rect 3869 8166 3921 8172
rect 4030 7086 4166 15920
rect 8408 14641 8460 14647
rect 8408 14583 8460 14589
rect 7297 14388 7989 14405
rect 7297 14205 7325 14388
rect 7956 14205 7989 14388
rect 7297 14189 7989 14205
rect 7759 13582 8167 13618
rect 7759 13312 7794 13582
rect 8130 13312 8167 13582
rect 7759 13275 8167 13312
rect 8416 12855 8452 14583
rect 8408 12849 8460 12855
rect 8408 12791 8460 12797
rect 8146 11719 8282 11759
rect 7548 11292 8282 11719
rect 7297 9755 7989 9772
rect 7297 9572 7325 9755
rect 7956 9572 7989 9755
rect 7297 9556 7989 9572
rect 7759 9089 8027 9125
rect 7759 8679 7794 9089
rect 7990 8679 8027 9089
rect 7759 8642 8027 8679
rect 4030 6654 4548 7086
rect 3870 5291 3922 5297
rect 3870 5233 3922 5239
rect 3878 3590 3914 5233
rect 3870 3584 3922 3590
rect 3870 3526 3922 3532
rect 3040 2021 3766 2453
rect 3630 1342 3766 2021
rect 4030 1342 4166 6654
rect 7297 5122 7989 5139
rect 7297 4939 7325 5122
rect 7956 4939 7989 5122
rect 7297 4923 7989 4939
rect 7759 4456 8027 4492
rect 7759 4046 7794 4456
rect 7990 4046 8027 4456
rect 7759 4009 8027 4046
rect 8146 2453 8282 11292
rect 8402 10008 8454 10014
rect 8402 9950 8454 9956
rect 8410 8224 8446 9950
rect 8402 8218 8454 8224
rect 8402 8160 8454 8166
rect 8546 7086 8682 15920
rect 12909 14725 12961 14731
rect 12909 14667 12961 14673
rect 11813 14388 12505 14405
rect 11813 14205 11841 14388
rect 12472 14205 12505 14388
rect 11813 14189 12505 14205
rect 12275 13582 12683 13618
rect 12275 13312 12310 13582
rect 12646 13312 12683 13582
rect 12275 13275 12683 13312
rect 12917 12868 12953 14667
rect 12909 12862 12961 12868
rect 12909 12804 12961 12810
rect 12662 11719 12798 11743
rect 12050 11287 12798 11719
rect 11813 9755 12505 9772
rect 11813 9572 11841 9755
rect 12472 9572 12505 9755
rect 11813 9556 12505 9572
rect 12275 9089 12543 9124
rect 12275 8679 12310 9089
rect 12506 8679 12543 9089
rect 12275 8642 12543 8679
rect 8546 6654 9032 7086
rect 8403 5375 8455 5381
rect 8403 5317 8455 5323
rect 8411 3599 8447 5317
rect 8403 3593 8455 3599
rect 8403 3535 8455 3541
rect 7566 2021 8282 2453
rect 8146 1342 8282 2021
rect 8546 1342 8682 6654
rect 11813 5122 12505 5139
rect 11813 4939 11841 5122
rect 12472 4939 12505 5122
rect 11813 4923 12505 4939
rect 12275 4456 12543 4492
rect 12275 4046 12310 4456
rect 12506 4046 12543 4456
rect 12275 4009 12543 4046
rect 12662 2453 12798 11287
rect 12920 10092 12972 10098
rect 12920 10034 12972 10040
rect 12928 8230 12964 10034
rect 12920 8224 12972 8230
rect 12920 8166 12972 8172
rect 13062 7086 13198 15920
rect 17407 14725 17459 14731
rect 17407 14667 17459 14673
rect 16329 14388 17021 14405
rect 16329 14205 16357 14388
rect 16988 14205 17021 14388
rect 16329 14189 17021 14205
rect 16791 13582 17199 13618
rect 16791 13312 16826 13582
rect 17162 13312 17199 13582
rect 16791 13275 17199 13312
rect 17415 12862 17451 14667
rect 17407 12856 17459 12862
rect 17407 12798 17459 12804
rect 17178 11719 17314 11751
rect 16586 11287 17314 11719
rect 16329 9755 17021 9772
rect 16329 9572 16357 9755
rect 16988 9572 17021 9755
rect 16329 9556 17021 9572
rect 16791 9089 17059 9125
rect 16791 8679 16826 9089
rect 17022 8679 17059 9089
rect 16791 8642 17059 8679
rect 13062 6654 13534 7086
rect 12900 5459 12952 5465
rect 12900 5401 12952 5407
rect 12908 3599 12944 5401
rect 12900 3593 12952 3599
rect 12900 3535 12952 3541
rect 12068 2021 12798 2453
rect 12662 1342 12798 2021
rect 13062 1342 13198 6654
rect 16329 5122 17021 5139
rect 16329 4939 16357 5122
rect 16988 4939 17021 5122
rect 16329 4923 17021 4939
rect 16791 4456 17059 4491
rect 16791 4046 16826 4456
rect 17022 4046 17059 4456
rect 16791 4009 17059 4046
rect 17178 2453 17314 11287
rect 17432 10092 17484 10098
rect 17432 10034 17484 10040
rect 17440 8233 17476 10034
rect 17432 8227 17484 8233
rect 17432 8169 17484 8175
rect 17578 7086 17714 15920
rect 21951 14641 22003 14647
rect 21951 14583 22003 14589
rect 20845 14388 21537 14405
rect 20845 14205 20873 14388
rect 21504 14205 21537 14388
rect 20845 14189 21537 14205
rect 21307 13582 21715 13618
rect 21307 13312 21342 13582
rect 21678 13312 21715 13582
rect 21307 13275 21715 13312
rect 21959 12863 21995 14583
rect 21951 12857 22003 12863
rect 21951 12799 22003 12805
rect 21694 11719 21830 11759
rect 21086 11287 21830 11719
rect 20845 9755 21537 9772
rect 20845 9572 20873 9755
rect 21504 9572 21537 9755
rect 20845 9556 21537 9572
rect 21307 9089 21575 9125
rect 21307 8679 21342 9089
rect 21538 8679 21575 9089
rect 21307 8642 21575 8679
rect 17578 6654 18060 7086
rect 17445 5459 17497 5465
rect 17445 5401 17497 5407
rect 17453 3591 17489 5401
rect 17445 3585 17497 3591
rect 17445 3527 17497 3533
rect 16604 2021 17314 2453
rect 17178 1342 17314 2021
rect 17578 1342 17714 6654
rect 20845 5122 21537 5139
rect 20845 4939 20873 5122
rect 21504 4939 21537 5122
rect 20845 4923 21537 4939
rect 21307 4456 21575 4492
rect 21307 4046 21342 4456
rect 21538 4046 21575 4456
rect 21307 4009 21575 4046
rect 21694 2453 21830 11287
rect 21944 10008 21996 10014
rect 21944 9950 21996 9956
rect 21952 8233 21988 9950
rect 21944 8227 21996 8233
rect 21944 8169 21996 8175
rect 22094 7086 22230 15920
rect 26495 14557 26547 14563
rect 26495 14499 26547 14505
rect 25361 14388 26053 14405
rect 25361 14205 25389 14388
rect 26020 14205 26053 14388
rect 25361 14189 26053 14205
rect 25823 13582 26231 13618
rect 25823 13312 25858 13582
rect 26194 13312 26231 13582
rect 25823 13275 26231 13312
rect 26503 12862 26539 14499
rect 26495 12856 26547 12862
rect 26495 12798 26547 12804
rect 26210 11719 26346 11759
rect 25614 11287 26346 11719
rect 25361 9755 26053 9772
rect 25361 9572 25389 9755
rect 26020 9572 26053 9755
rect 25361 9556 26053 9572
rect 25823 9089 26091 9125
rect 25823 8679 25858 9089
rect 26054 8679 26091 9089
rect 25823 8642 26091 8679
rect 22094 6654 22578 7086
rect 21958 5375 22010 5381
rect 21958 5317 22010 5323
rect 21966 3591 22002 5317
rect 21958 3585 22010 3591
rect 21958 3527 22010 3533
rect 21104 2021 21830 2453
rect 21694 1342 21830 2021
rect 22094 1342 22230 6654
rect 25361 5122 26053 5139
rect 25361 4939 25389 5122
rect 26020 4939 26053 5122
rect 25361 4923 26053 4939
rect 25823 4456 26091 4492
rect 25823 4046 25858 4456
rect 26054 4046 26091 4456
rect 25823 4009 26091 4046
rect 26210 2453 26346 11287
rect 26409 10097 26461 10103
rect 26409 10039 26461 10045
rect 26417 8230 26453 10039
rect 26507 9939 26559 9945
rect 26507 9881 26559 9887
rect 26409 8224 26461 8230
rect 26409 8166 26461 8172
rect 26515 5465 26551 9881
rect 29877 9755 30569 9772
rect 29877 9572 29905 9755
rect 30536 9572 30569 9755
rect 29877 9556 30569 9572
rect 30339 8949 30747 8985
rect 30339 8679 30374 8949
rect 30710 8679 30747 8949
rect 30339 8642 30747 8679
rect 30930 8224 30982 8230
rect 30930 8166 30982 8172
rect 26610 7086 26746 7096
rect 26610 6654 27080 7086
rect 26507 5459 26559 5465
rect 26507 5401 26559 5407
rect 26421 5291 26473 5297
rect 26421 5233 26473 5239
rect 26429 3601 26465 5233
rect 26421 3595 26473 3601
rect 26421 3537 26473 3543
rect 25622 2021 26346 2453
rect 26210 1342 26346 2021
rect 26610 1342 26746 6654
rect 29877 5122 30569 5139
rect 29877 4939 29905 5122
rect 30536 4939 30569 5122
rect 29877 4923 30569 4939
rect 30339 4316 30747 4352
rect 30339 4046 30374 4316
rect 30710 4046 30747 4316
rect 30339 4009 30747 4046
rect 30726 2453 30862 2484
rect 30132 2021 30862 2453
rect 30726 1342 30862 2021
rect 30938 770 30974 8166
rect 31025 5375 31061 9943
rect 34393 9755 35085 9772
rect 34393 9572 34421 9755
rect 35052 9572 35085 9755
rect 34393 9556 35085 9572
rect 34855 8949 35263 8985
rect 34855 8679 34890 8949
rect 35226 8679 35263 8949
rect 34855 8642 35263 8679
rect 35441 8237 35493 8243
rect 35441 8179 35493 8185
rect 31126 7086 31262 7121
rect 31126 6654 31606 7086
rect 31011 5323 31017 5375
rect 31069 5323 31075 5375
rect 31126 1342 31262 6654
rect 34393 5122 35085 5139
rect 34393 4939 34421 5122
rect 35052 4939 35085 5122
rect 34393 4923 35085 4939
rect 34855 4316 35263 4352
rect 34855 4046 34890 4316
rect 35226 4046 35263 4316
rect 34855 4009 35263 4046
rect 35242 2453 35378 2503
rect 34660 2021 35378 2453
rect 35242 1342 35378 2021
rect 30930 764 30982 770
rect 30930 706 30982 712
rect 35449 597 35485 8179
rect 35553 5297 35589 9939
rect 38909 9755 39602 9772
rect 38909 9572 38937 9755
rect 39568 9572 39602 9755
rect 38909 9556 39602 9572
rect 39371 9089 39639 9125
rect 39371 8679 39406 9089
rect 39602 8679 39639 9089
rect 39371 8642 39639 8679
rect 39681 8239 39709 9932
rect 39669 8233 39721 8239
rect 39669 8175 39721 8181
rect 35642 7086 35778 7130
rect 35642 6654 36126 7086
rect 35545 5291 35597 5297
rect 35545 5233 35597 5239
rect 35642 1342 35778 6654
rect 38909 5122 39601 5139
rect 38909 4939 38937 5122
rect 39568 4939 39601 5122
rect 38909 4923 39601 4939
rect 39371 4316 39779 4352
rect 39371 4046 39406 4316
rect 39742 4046 39779 4316
rect 39371 4009 39779 4046
rect 39982 3598 40010 9952
rect 39973 3592 40025 3598
rect 39973 3534 40025 3540
rect 40066 3309 40094 9952
rect 40400 7941 40428 9924
rect 43425 9755 44117 9772
rect 43425 9572 43453 9755
rect 44084 9572 44117 9755
rect 43425 9556 44117 9572
rect 43887 9089 44155 9125
rect 43887 8679 43922 9089
rect 44118 8679 44155 9089
rect 43887 8642 44155 8679
rect 40388 7935 40440 7941
rect 40388 7877 40440 7883
rect 40158 7086 40294 7092
rect 40158 6654 40626 7086
rect 40051 3303 40103 3309
rect 40051 3245 40103 3251
rect 39758 2453 39894 2484
rect 39170 2021 39894 2453
rect 39758 1342 39894 2021
rect 40158 1342 40294 6654
rect 43425 5122 44117 5139
rect 43425 4939 43453 5122
rect 44084 4939 44117 5122
rect 43425 4923 44117 4939
rect 43887 4456 44155 4492
rect 43887 4046 43922 4456
rect 44118 4046 44155 4456
rect 43887 4009 44155 4046
rect 44274 2453 44410 2503
rect 43680 2021 44410 2453
rect 44274 1342 44410 2021
rect 35441 591 35493 597
rect 35441 533 35493 539
<< via2 >>
rect 2809 18838 3440 19021
rect 3278 17945 3614 18215
rect 7325 18838 7956 19021
rect 7794 17945 8130 18215
rect 11841 18838 12472 19021
rect 12310 17945 12646 18215
rect 16357 18838 16988 19021
rect 16826 17945 17162 18215
rect 20873 18838 21504 19021
rect 21342 17945 21678 18215
rect 25389 18838 26020 19021
rect 25858 17945 26194 18215
rect 631 16514 2857 16663
rect 5147 16514 7373 16663
rect 9663 16514 11889 16663
rect 14179 16514 16405 16663
rect 18695 16514 20921 16663
rect 23211 16514 25437 16663
rect 499 15060 2830 15172
rect 2809 14205 3440 14388
rect 3278 13312 3614 13582
rect 631 11881 2857 12030
rect 499 10427 2830 10539
rect 2809 9572 3440 9755
rect 3278 8679 3474 9089
rect 631 7248 2857 7397
rect 499 5794 2830 5906
rect 2809 4939 3440 5122
rect 3278 4046 3474 4456
rect 631 2615 2857 2764
rect 5015 15060 7346 15172
rect 7325 14205 7956 14388
rect 7794 13312 8130 13582
rect 5147 11881 7373 12030
rect 5015 10427 7346 10539
rect 7325 9572 7956 9755
rect 7794 8679 7990 9089
rect 5147 7248 7373 7397
rect 5015 5794 7346 5906
rect 7325 4939 7956 5122
rect 7794 4046 7990 4456
rect 5147 2615 7373 2764
rect 9531 15060 11862 15172
rect 11841 14205 12472 14388
rect 12310 13312 12646 13582
rect 9663 11881 11889 12030
rect 9531 10427 11862 10539
rect 11841 9572 12472 9755
rect 12310 8679 12506 9089
rect 9663 7248 11889 7397
rect 9531 5794 11862 5906
rect 11841 4939 12472 5122
rect 12310 4046 12506 4456
rect 9663 2615 11889 2764
rect 14047 15060 16378 15172
rect 16357 14205 16988 14388
rect 16826 13312 17162 13582
rect 14179 11881 16405 12030
rect 14047 10427 16378 10539
rect 16357 9572 16988 9755
rect 16826 8679 17022 9089
rect 14179 7248 16405 7397
rect 14047 5794 16378 5906
rect 16357 4939 16988 5122
rect 16826 4046 17022 4456
rect 14179 2615 16405 2764
rect 18563 15060 20894 15172
rect 20873 14205 21504 14388
rect 21342 13312 21678 13582
rect 18695 11881 20921 12030
rect 18563 10427 20894 10539
rect 20873 9572 21504 9755
rect 21342 8679 21538 9089
rect 18695 7248 20921 7397
rect 18563 5794 20894 5906
rect 20873 4939 21504 5122
rect 21342 4046 21538 4456
rect 18695 2615 20921 2764
rect 23079 15060 25410 15172
rect 25389 14205 26020 14388
rect 25858 13312 26194 13582
rect 23211 11881 25437 12030
rect 23079 10427 25410 10539
rect 25389 9572 26020 9755
rect 25858 8679 26054 9089
rect 23211 7248 25437 7397
rect 23079 5794 25410 5906
rect 25389 4939 26020 5122
rect 25858 4046 26054 4456
rect 23211 2615 25437 2764
rect 29905 9572 30536 9755
rect 30374 8679 30710 8949
rect 27727 7248 29953 7397
rect 27595 5794 29926 5906
rect 29905 4939 30536 5122
rect 30374 4046 30710 4316
rect 27727 2615 29953 2764
rect 499 1161 2830 1273
rect 5015 1161 7346 1273
rect 9531 1161 11862 1273
rect 14047 1161 16378 1273
rect 18563 1161 20894 1273
rect 23079 1161 25410 1273
rect 27595 1161 29926 1273
rect 34421 9572 35052 9755
rect 34890 8679 35226 8949
rect 32243 7248 34469 7397
rect 32111 5794 34442 5906
rect 34421 4939 35052 5122
rect 34890 4046 35226 4316
rect 32243 2615 34469 2764
rect 32111 1161 34442 1273
rect 38937 9572 39568 9755
rect 39406 8679 39602 9089
rect 36759 7248 38985 7397
rect 36627 5794 38958 5906
rect 38937 4939 39568 5122
rect 39406 4046 39742 4316
rect 43453 9572 44084 9755
rect 43922 8679 44118 9089
rect 41275 7248 43501 7397
rect 36759 2615 38985 2764
rect 41143 5794 43474 5906
rect 43453 4939 44084 5122
rect 43922 4046 44118 4456
rect 41275 2615 43501 2764
rect 36627 1161 38958 1273
rect 41143 1161 43474 1273
<< metal3 >>
rect -935 19036 26452 19053
rect -935 19021 8160 19036
rect -935 18838 2809 19021
rect 3440 18838 7325 19021
rect 7956 18838 8160 19021
rect -935 18837 8160 18838
rect 8618 19021 26452 19036
rect 8618 18838 11841 19021
rect 12472 18838 16357 19021
rect 16988 18838 20873 19021
rect 21504 18838 25389 19021
rect 26020 18838 26452 19021
rect 8618 18837 26452 18838
rect -935 18826 26452 18837
rect 2781 18822 3473 18826
rect 7297 18822 7989 18826
rect 11813 18822 12505 18826
rect 16329 18822 17021 18826
rect 20845 18822 21537 18826
rect 25361 18822 26053 18826
rect 40 18245 26459 18259
rect 40 18215 12743 18245
rect 40 18083 3278 18215
rect 3243 17945 3278 18083
rect 3614 18083 7794 18215
rect 3614 17945 3651 18083
rect 3243 17908 3651 17945
rect 7759 17945 7794 18083
rect 8130 18083 12310 18215
rect 8130 17945 8167 18083
rect 7759 17908 8167 17945
rect 12275 17945 12310 18083
rect 12646 18097 12743 18215
rect 13150 18215 26459 18245
rect 13150 18097 16826 18215
rect 12646 18083 16826 18097
rect 12646 17945 12683 18083
rect 12275 17908 12683 17945
rect 16791 17945 16826 18083
rect 17162 18083 21342 18215
rect 17162 17945 17199 18083
rect 16791 17908 17199 17945
rect 21307 17945 21342 18083
rect 21678 18083 25858 18215
rect 21678 17945 21715 18083
rect 21307 17908 21715 17945
rect 25823 17945 25858 18083
rect 26194 18083 26459 18215
rect 26194 17945 26231 18083
rect 25823 17908 26231 17945
rect -111 16683 26308 16688
rect -111 16678 26393 16683
rect -111 16663 3658 16678
rect -111 16514 631 16663
rect 2857 16517 3658 16663
rect 4123 16668 26393 16678
rect 4123 16663 21715 16668
rect 4123 16517 5147 16663
rect 2857 16514 5147 16517
rect 7373 16514 9663 16663
rect 11889 16514 14179 16663
rect 16405 16514 18695 16663
rect 20921 16520 21715 16663
rect 22173 16663 26393 16668
rect 22173 16520 23211 16663
rect 20921 16514 23211 16520
rect 25437 16514 26393 16663
rect -111 16512 26393 16514
rect -26 16507 26393 16512
rect 469 16500 2955 16507
rect 4985 16500 7471 16507
rect 9501 16500 11987 16507
rect 14017 16500 16503 16507
rect 18533 16500 21019 16507
rect 23049 16500 25535 16507
rect -756 15360 25864 15792
rect 377 15188 2938 15209
rect 4893 15188 7454 15209
rect 9409 15188 11970 15209
rect 13925 15188 16486 15209
rect 18441 15188 21002 15209
rect 22957 15188 25518 15209
rect -929 15180 26372 15188
rect -929 15019 -894 15180
rect -429 15172 26372 15180
rect -429 15060 499 15172
rect 2830 15060 5015 15172
rect 7346 15060 9531 15172
rect 11862 15060 14047 15172
rect 16378 15060 17226 15172
rect -429 15024 17226 15060
rect 17684 15060 18563 15172
rect 20894 15060 23079 15172
rect 25410 15060 26372 15172
rect 17684 15024 26372 15060
rect -429 15019 26372 15024
rect -929 15012 26372 15019
rect -930 14407 26452 14420
rect -930 14388 8164 14407
rect -930 14205 2809 14388
rect 3440 14205 7325 14388
rect 7956 14208 8164 14388
rect 8622 14388 26452 14407
rect 8622 14208 11841 14388
rect 7956 14205 11841 14208
rect 12472 14205 16357 14388
rect 16988 14205 20873 14388
rect 21504 14205 25389 14388
rect 26020 14205 26452 14388
rect -930 14193 26452 14205
rect 2781 14189 3473 14193
rect 7297 14189 7989 14193
rect 11813 14189 12505 14193
rect 16329 14189 17021 14193
rect 20845 14189 21537 14193
rect 25361 14189 26053 14193
rect 40 13609 26459 13626
rect 40 13582 12734 13609
rect 40 13450 3278 13582
rect 3243 13312 3278 13450
rect 3614 13450 7794 13582
rect 3614 13312 3651 13450
rect 3243 13275 3651 13312
rect 7759 13312 7794 13450
rect 8130 13450 12310 13582
rect 8130 13312 8167 13450
rect 7759 13275 8167 13312
rect 12275 13312 12310 13450
rect 12646 13461 12734 13582
rect 13152 13582 26459 13609
rect 13152 13461 16826 13582
rect 12646 13450 16826 13461
rect 12646 13312 12683 13450
rect 12275 13275 12683 13312
rect 16791 13312 16826 13450
rect 17162 13450 21342 13582
rect 17162 13312 17199 13450
rect 16791 13275 17199 13312
rect 21307 13312 21342 13450
rect 21678 13450 25858 13582
rect 21678 13312 21715 13450
rect 21307 13275 21715 13312
rect 25823 13312 25858 13450
rect 26194 13450 26459 13582
rect 26194 13312 26231 13450
rect 25823 13275 26231 13312
rect 469 12050 2955 12053
rect 4985 12050 7471 12053
rect 9501 12050 11987 12053
rect 14017 12050 16503 12053
rect 18533 12050 21019 12053
rect 23049 12050 25535 12053
rect -26 12044 26393 12050
rect -26 12030 3658 12044
rect -26 11881 631 12030
rect 2857 11883 3658 12030
rect 4123 12036 26393 12044
rect 4123 12030 21719 12036
rect 4123 11883 5147 12030
rect 2857 11881 5147 11883
rect 7373 11881 9663 12030
rect 11889 11881 14179 12030
rect 16405 11881 18695 12030
rect 20921 11888 21719 12030
rect 22177 12030 26393 12036
rect 22177 11888 23211 12030
rect 20921 11881 23211 11888
rect 25437 11881 26393 12030
rect -26 11874 26393 11881
rect 469 11867 2955 11874
rect 4985 11867 7471 11874
rect 9501 11867 11987 11874
rect 14017 11867 16503 11874
rect 18533 11867 21019 11874
rect 23049 11867 25535 11874
rect -790 10727 25864 11159
rect 377 10555 2938 10576
rect 4893 10555 7454 10576
rect 9409 10555 11970 10576
rect 13925 10555 16486 10576
rect 18441 10555 21002 10576
rect 22957 10555 25518 10576
rect -909 10551 26372 10555
rect -909 10390 -894 10551
rect -429 10539 26372 10551
rect -429 10427 499 10539
rect 2830 10427 5015 10539
rect 7346 10427 9531 10539
rect 11862 10427 14047 10539
rect 16378 10536 18563 10539
rect 16378 10427 17224 10536
rect -429 10390 17224 10427
rect -909 10388 17224 10390
rect 17682 10427 18563 10536
rect 20894 10427 23079 10539
rect 25410 10427 26372 10539
rect 17682 10388 26372 10427
rect -909 10379 26372 10388
rect -910 9773 44089 9787
rect -910 9755 8164 9773
rect -910 9572 2809 9755
rect 3440 9572 7325 9755
rect 7956 9572 8164 9755
rect 8626 9772 44089 9773
rect 8626 9755 44117 9772
rect 8626 9572 11841 9755
rect 12472 9572 16357 9755
rect 16988 9572 20873 9755
rect 21504 9572 25389 9755
rect 26020 9572 29905 9755
rect 30536 9572 34421 9755
rect 35052 9572 38937 9755
rect 39568 9572 43453 9755
rect 44084 9572 44117 9755
rect -910 9560 44117 9572
rect 2781 9555 3473 9560
rect 7297 9556 7989 9560
rect 11813 9556 12505 9560
rect 16329 9556 17021 9560
rect 20845 9556 21537 9560
rect 25361 9556 26053 9560
rect 29877 9556 30569 9560
rect 34393 9556 35085 9560
rect 38909 9556 39601 9560
rect 43425 9556 44117 9560
rect 3243 9089 3512 9125
rect 3243 8993 3278 9089
rect 40 8817 3278 8993
rect 3243 8679 3278 8817
rect 3474 8993 3512 9089
rect 7758 9089 8027 9125
rect 7758 8993 7794 9089
rect 3474 8817 7794 8993
rect 3474 8679 3511 8817
rect 3243 8642 3511 8679
rect 7759 8679 7794 8817
rect 7990 8993 8027 9089
rect 12275 9089 12544 9124
rect 12275 8993 12310 9089
rect 7990 8817 12310 8993
rect 7990 8679 8027 8817
rect 7759 8642 8027 8679
rect 12275 8679 12310 8817
rect 12506 8993 12544 9089
rect 16791 9089 17059 9125
rect 16791 8993 16826 9089
rect 12506 8982 16826 8993
rect 12506 8834 12690 8982
rect 13148 8834 16826 8982
rect 12506 8817 16826 8834
rect 12506 8679 12543 8817
rect 12275 8642 12543 8679
rect 16791 8679 16826 8817
rect 17022 8993 17059 9089
rect 21307 9089 21575 9125
rect 21307 8993 21342 9089
rect 17022 8817 21342 8993
rect 17022 8679 17059 8817
rect 16791 8642 17059 8679
rect 21307 8679 21342 8817
rect 21538 8993 21575 9089
rect 25823 9089 26091 9125
rect 25823 8993 25858 9089
rect 21538 8817 25858 8993
rect 21538 8679 21575 8817
rect 21307 8642 21575 8679
rect 25823 8679 25858 8817
rect 26054 8993 26091 9089
rect 39371 9089 39639 9125
rect 39371 8993 39406 9089
rect 26054 8949 39406 8993
rect 26054 8817 30374 8949
rect 26054 8679 26091 8817
rect 25823 8642 26091 8679
rect 30339 8679 30374 8817
rect 30710 8817 34890 8949
rect 30710 8679 30747 8817
rect 30339 8642 30747 8679
rect 34855 8679 34890 8817
rect 35226 8817 39406 8949
rect 35226 8679 35263 8817
rect 34855 8642 35263 8679
rect 39371 8679 39406 8817
rect 39602 8993 39639 9089
rect 43887 9089 44155 9125
rect 43887 8993 43922 9089
rect 39602 8817 43922 8993
rect 39602 8679 39639 8817
rect 39371 8642 39639 8679
rect 43887 8679 43922 8817
rect 44118 8993 44155 9089
rect 44118 8817 44179 8993
rect 44118 8679 44155 8817
rect 43887 8642 44155 8679
rect 469 7417 2955 7420
rect 4985 7417 7471 7420
rect 9501 7417 11987 7420
rect 14017 7417 16503 7420
rect 18533 7417 21019 7420
rect 23049 7417 25535 7420
rect 27565 7417 30051 7420
rect 32081 7417 34567 7420
rect 36597 7417 39083 7420
rect 41113 7417 43599 7420
rect -26 7413 44096 7417
rect -26 7397 3656 7413
rect -26 7248 631 7397
rect 2857 7252 3656 7397
rect 4121 7403 44096 7413
rect 4121 7397 21715 7403
rect 4121 7252 5147 7397
rect 2857 7248 5147 7252
rect 7373 7248 9663 7397
rect 11889 7248 14179 7397
rect 16405 7248 18695 7397
rect 20921 7255 21715 7397
rect 22173 7397 44096 7403
rect 22173 7255 23211 7397
rect 20921 7248 23211 7255
rect 25437 7248 27727 7397
rect 29953 7248 32243 7397
rect 34469 7248 36759 7397
rect 38985 7248 41275 7397
rect 43501 7248 44096 7397
rect -26 7241 44096 7248
rect 469 7234 2955 7241
rect 4985 7234 7471 7241
rect 9501 7234 11987 7241
rect 14017 7234 16503 7241
rect 18533 7234 21019 7241
rect 23049 7234 25535 7241
rect 27565 7234 30051 7241
rect 32081 7234 34567 7241
rect 36597 7234 39083 7241
rect 41113 7234 43599 7241
rect -670 6094 43778 6526
rect 377 5922 2938 5943
rect 4893 5922 7454 5943
rect 9409 5922 11970 5943
rect 13925 5922 16486 5943
rect 18441 5922 21002 5943
rect 22957 5922 25518 5943
rect 27473 5922 30034 5943
rect 31989 5922 34550 5943
rect 36505 5922 39066 5943
rect 41021 5922 43582 5943
rect -909 5914 44179 5922
rect -909 5753 -892 5914
rect -427 5909 44179 5914
rect -427 5906 17228 5909
rect -427 5794 499 5906
rect 2830 5794 5015 5906
rect 7346 5794 9531 5906
rect 11862 5794 14047 5906
rect 16378 5794 17228 5906
rect -427 5761 17228 5794
rect 17686 5906 44179 5909
rect 17686 5794 18563 5906
rect 20894 5794 23079 5906
rect 25410 5794 27595 5906
rect 29926 5794 32111 5906
rect 34442 5794 36627 5906
rect 38958 5794 41143 5906
rect 43474 5794 44179 5906
rect 17686 5761 44179 5794
rect -427 5753 44179 5761
rect -909 5746 44179 5753
rect -930 5142 44161 5154
rect -930 5122 8162 5142
rect -930 4939 2809 5122
rect 3440 4939 7325 5122
rect 7956 4941 8162 5122
rect 8624 5122 44161 5142
rect 8624 4941 11841 5122
rect 7956 4939 11841 4941
rect 12472 4939 16357 5122
rect 16988 4939 20873 5122
rect 21504 4939 25389 5122
rect 26020 4939 29905 5122
rect 30536 4939 34421 5122
rect 35052 4939 38937 5122
rect 39568 4939 43453 5122
rect 44084 4939 44161 5122
rect -930 4927 44161 4939
rect 2781 4923 3473 4927
rect 7297 4923 7989 4927
rect 11813 4923 12505 4927
rect 16329 4923 17021 4927
rect 20845 4923 21537 4927
rect 25361 4923 26053 4927
rect 29877 4923 30569 4927
rect 34393 4923 35085 4927
rect 38909 4923 39601 4927
rect 43425 4923 44117 4927
rect 3243 4456 3511 4492
rect 3243 4360 3278 4456
rect 40 4184 3278 4360
rect 3243 4046 3278 4184
rect 3474 4360 3511 4456
rect 7759 4456 8027 4492
rect 7759 4360 7794 4456
rect 3474 4184 7794 4360
rect 3474 4046 3511 4184
rect 3243 4009 3511 4046
rect 7759 4046 7794 4184
rect 7990 4360 8027 4456
rect 12275 4456 12543 4492
rect 12275 4360 12310 4456
rect 7990 4184 12310 4360
rect 7990 4046 8027 4184
rect 7759 4009 8027 4046
rect 12275 4046 12310 4184
rect 12506 4360 12543 4456
rect 16791 4456 17059 4491
rect 16791 4360 16826 4456
rect 12506 4342 16826 4360
rect 12506 4194 12692 4342
rect 13150 4194 16826 4342
rect 12506 4184 16826 4194
rect 12506 4046 12543 4184
rect 12275 4009 12543 4046
rect 16791 4046 16826 4184
rect 17022 4360 17059 4456
rect 21307 4456 21575 4492
rect 21307 4360 21342 4456
rect 17022 4184 21342 4360
rect 17022 4046 17059 4184
rect 16791 4009 17059 4046
rect 21307 4046 21342 4184
rect 21538 4360 21575 4456
rect 25823 4456 26091 4492
rect 25823 4360 25858 4456
rect 21538 4184 25858 4360
rect 21538 4046 21575 4184
rect 21307 4009 21575 4046
rect 25823 4046 25858 4184
rect 26054 4360 26091 4456
rect 43887 4456 44155 4492
rect 43887 4360 43922 4456
rect 26054 4316 43922 4360
rect 26054 4184 30374 4316
rect 26054 4046 26091 4184
rect 25823 4009 26091 4046
rect 30339 4046 30374 4184
rect 30710 4184 34890 4316
rect 30710 4046 30747 4184
rect 30339 4009 30747 4046
rect 34855 4046 34890 4184
rect 35226 4184 39406 4316
rect 35226 4046 35263 4184
rect 34855 4009 35263 4046
rect 39371 4046 39406 4184
rect 39742 4184 43922 4316
rect 39742 4046 39779 4184
rect 39371 4009 39779 4046
rect 43887 4046 43922 4184
rect 44118 4360 44155 4456
rect 44118 4184 44210 4360
rect 44118 4046 44155 4184
rect 43887 4009 44155 4046
rect 469 2784 2955 2787
rect 4985 2784 7471 2787
rect 9501 2784 11987 2787
rect 14017 2784 16503 2787
rect 18533 2784 21019 2787
rect 23049 2784 25535 2787
rect 27565 2784 30051 2787
rect 32081 2784 34567 2787
rect 36597 2784 39083 2787
rect 41113 2784 43599 2787
rect -26 2778 44096 2784
rect -26 2764 3658 2778
rect -26 2615 631 2764
rect 2857 2617 3658 2764
rect 4123 2767 44096 2778
rect 4123 2764 21715 2767
rect 4123 2617 5147 2764
rect 2857 2615 5147 2617
rect 7373 2615 9663 2764
rect 11889 2615 14179 2764
rect 16405 2615 18695 2764
rect 20921 2619 21715 2764
rect 22173 2764 44096 2767
rect 22173 2619 23211 2764
rect 20921 2615 23211 2619
rect 25437 2615 27727 2764
rect 29953 2615 32243 2764
rect 34469 2615 36759 2764
rect 38985 2615 41275 2764
rect 43501 2615 44096 2764
rect -26 2608 44096 2615
rect 469 2601 2955 2608
rect 4985 2601 7471 2608
rect 9501 2601 11987 2608
rect 14017 2601 16503 2608
rect 18533 2601 21019 2608
rect 23049 2601 25535 2608
rect 27565 2601 30051 2608
rect 32081 2601 34567 2608
rect 36597 2601 39083 2608
rect 41113 2601 43599 2608
rect -602 1461 43778 1893
rect 377 1289 2938 1310
rect 4893 1289 7454 1310
rect 9409 1289 11970 1310
rect 13925 1289 16486 1310
rect 18441 1289 21002 1310
rect 22957 1289 25518 1310
rect 27473 1289 30034 1310
rect 31989 1289 34550 1310
rect 36505 1289 39066 1310
rect 41021 1289 43582 1310
rect -929 1282 44085 1289
rect -929 1121 -894 1282
rect -429 1273 44085 1282
rect -429 1161 499 1273
rect 2830 1161 5015 1273
rect 7346 1161 9531 1273
rect 11862 1161 14047 1273
rect 16378 1272 18563 1273
rect 16378 1161 17226 1272
rect -429 1124 17226 1161
rect 17684 1161 18563 1272
rect 20894 1161 23079 1273
rect 25410 1161 27595 1273
rect 29926 1161 32111 1273
rect 34442 1161 36627 1273
rect 38958 1161 41143 1273
rect 43474 1161 44085 1273
rect 17684 1124 44085 1161
rect -429 1121 44085 1124
rect -929 1113 44085 1121
<< via3 >>
rect 8160 18837 8618 19036
rect 12743 18097 13150 18245
rect 3658 16517 4123 16678
rect 21715 16520 22173 16668
rect -894 15019 -429 15180
rect 17226 15024 17684 15172
rect 8164 14208 8622 14407
rect 12734 13461 13152 13609
rect 3658 11883 4123 12044
rect 21719 11888 22177 12036
rect -894 10390 -429 10551
rect 17224 10388 17682 10536
rect 8164 9572 8626 9773
rect 12690 8834 13148 8982
rect 3656 7252 4121 7413
rect 21715 7255 22173 7403
rect -892 5753 -427 5914
rect 17228 5761 17686 5909
rect 8162 4941 8624 5142
rect 12692 4194 13150 4342
rect 3658 2617 4123 2778
rect 21715 2619 22173 2767
rect -894 1121 -429 1282
rect 17226 1124 17684 1272
<< metal4 >>
rect -901 15180 -419 19102
rect -901 15019 -894 15180
rect -429 15019 -419 15180
rect -901 10551 -419 15019
rect -901 10390 -894 10551
rect -429 10390 -419 10551
rect -901 5914 -419 10390
rect -901 5753 -892 5914
rect -427 5753 -419 5914
rect -901 1282 -419 5753
rect -901 1121 -894 1282
rect -429 1121 -419 1282
rect -901 397 -419 1121
rect 3647 16678 4129 19102
rect 3647 16517 3658 16678
rect 4123 16517 4129 16678
rect 3647 12044 4129 16517
rect 3647 11883 3658 12044
rect 4123 11883 4129 12044
rect 3647 7413 4129 11883
rect 3647 7252 3656 7413
rect 4121 7252 4129 7413
rect 3647 2778 4129 7252
rect 3647 2617 3658 2778
rect 4123 2617 4129 2778
rect 3647 397 4129 2617
rect 8151 19036 8633 19102
rect 8151 18837 8160 19036
rect 8618 18837 8633 19036
rect 8151 14407 8633 18837
rect 8151 14208 8164 14407
rect 8622 14208 8633 14407
rect 8151 9773 8633 14208
rect 8151 9572 8164 9773
rect 8626 9572 8633 9773
rect 8151 5142 8633 9572
rect 8151 4941 8162 5142
rect 8624 4941 8633 5142
rect 8151 397 8633 4941
rect 12679 18245 13161 19118
rect 12679 18097 12743 18245
rect 13150 18097 13161 18245
rect 12679 13609 13161 18097
rect 12679 13461 12734 13609
rect 13152 13461 13161 13609
rect 12679 8982 13161 13461
rect 12679 8834 12690 8982
rect 13148 8834 13161 8982
rect 12679 4342 13161 8834
rect 12679 4194 12692 4342
rect 13150 4194 13161 4342
rect 12679 413 13161 4194
rect 17214 15172 17696 19102
rect 17214 15024 17226 15172
rect 17684 15024 17696 15172
rect 17214 10536 17696 15024
rect 17214 10388 17224 10536
rect 17682 10388 17696 10536
rect 17214 5909 17696 10388
rect 17214 5761 17228 5909
rect 17686 5761 17696 5909
rect 17214 1272 17696 5761
rect 17214 1124 17226 1272
rect 17684 1124 17696 1272
rect 17214 397 17696 1124
rect 21700 16668 22182 19102
rect 21700 16520 21715 16668
rect 22173 16520 22182 16668
rect 21700 12036 22182 16520
rect 21700 11888 21719 12036
rect 22177 11888 22182 12036
rect 21700 7403 22182 11888
rect 21700 7255 21715 7403
rect 22173 7255 22182 7403
rect 21700 2767 22182 7255
rect 21700 2619 21715 2767
rect 22173 2619 22182 2767
rect 21700 397 22182 2619
use cv3_via2_36cut  cv3_via2_36cut_0
timestamp 1719173892
transform 1 0 -550582 0 1 -90682
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_1
timestamp 1719173892
transform 1 0 -548960 0 1 -90678
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_2
timestamp 1719173892
transform 1 0 -553476 0 1 -90678
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_3
timestamp 1719173892
transform 1 0 -555098 0 1 -90682
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_4
timestamp 1719173892
transform 1 0 -546066 0 1 -90682
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_5
timestamp 1719173892
transform 1 0 -544444 0 1 -90678
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_6
timestamp 1719173892
transform 1 0 -541550 0 1 -90682
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_7
timestamp 1719173892
transform 1 0 -539928 0 1 -90678
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_8
timestamp 1719173892
transform 1 0 -537034 0 1 -90682
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_9
timestamp 1719173892
transform 1 0 -535412 0 1 -90678
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_10
timestamp 1719173892
transform 1 0 -532518 0 1 -90682
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_11
timestamp 1719173892
transform 1 0 -530896 0 1 -90678
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_12
timestamp 1719173892
transform 1 0 -528002 0 1 -90682
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_13
timestamp 1719173892
transform 1 0 -526380 0 1 -90678
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_14
timestamp 1719173892
transform 1 0 -523486 0 1 -90682
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_15
timestamp 1719173892
transform 1 0 -521864 0 1 -90678
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_16
timestamp 1719173892
transform 1 0 -518970 0 1 -90682
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_17
timestamp 1719173892
transform 1 0 -517348 0 1 -90678
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_18
timestamp 1719173892
transform 1 0 -555098 0 1 -86049
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_19
timestamp 1719173892
transform 1 0 -553476 0 1 -86045
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_20
timestamp 1719173892
transform 1 0 -514454 0 1 -90682
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_21
timestamp 1719173892
transform 1 0 -512832 0 1 -90678
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_22
timestamp 1719173892
transform 1 0 -514454 0 1 -86049
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_23
timestamp 1719173892
transform 1 0 -512832 0 1 -86045
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_24
timestamp 1719173892
transform 1 0 -518970 0 1 -86049
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_25
timestamp 1719173892
transform 1 0 -517348 0 1 -86045
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_26
timestamp 1719173892
transform 1 0 -523486 0 1 -86049
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_27
timestamp 1719173892
transform 1 0 -521864 0 1 -86045
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_28
timestamp 1719173892
transform 1 0 -526380 0 1 -86045
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_29
timestamp 1719173892
transform 1 0 -528002 0 1 -86049
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_30
timestamp 1719173892
transform 1 0 -532518 0 1 -86049
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_31
timestamp 1719173892
transform 1 0 -530896 0 1 -86045
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_32
timestamp 1719173892
transform 1 0 -537034 0 1 -86049
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_33
timestamp 1719173892
transform 1 0 -535412 0 1 -86045
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_34
timestamp 1719173892
transform 1 0 -541550 0 1 -86049
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_35
timestamp 1719173892
transform 1 0 -539928 0 1 -86045
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_36
timestamp 1719173892
transform 1 0 -546066 0 1 -86049
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_37
timestamp 1719173892
transform 1 0 -544444 0 1 -86045
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_38
timestamp 1719173892
transform 1 0 -550582 0 1 -86049
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_39
timestamp 1719173892
transform 1 0 -548960 0 1 -86045
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_40
timestamp 1719173892
transform 1 0 -532518 0 1 -81416
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_41
timestamp 1719173892
transform 1 0 -530896 0 1 -81412
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_42
timestamp 1719173892
transform 1 0 -555098 0 1 -81416
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_43
timestamp 1719173892
transform 1 0 -553476 0 1 -81412
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_44
timestamp 1719173892
transform 1 0 -550582 0 1 -81416
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_45
timestamp 1719173892
transform 1 0 -548960 0 1 -81412
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_46
timestamp 1719173892
transform 1 0 -546066 0 1 -81416
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_47
timestamp 1719173892
transform 1 0 -544444 0 1 -81412
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_48
timestamp 1719173892
transform 1 0 -541550 0 1 -81416
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_49
timestamp 1719173892
transform 1 0 -539928 0 1 -81412
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_50
timestamp 1719173892
transform 1 0 -537034 0 1 -81416
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_51
timestamp 1719173892
transform 1 0 -535412 0 1 -81412
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_52
timestamp 1719173892
transform 1 0 -555098 0 1 -76783
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_53
timestamp 1719173892
transform 1 0 -553476 0 1 -76779
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_54
timestamp 1719173892
transform 1 0 -532518 0 1 -76783
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_55
timestamp 1719173892
transform 1 0 -530896 0 1 -76779
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_56
timestamp 1719173892
transform 1 0 -537034 0 1 -76783
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_57
timestamp 1719173892
transform 1 0 -535412 0 1 -76779
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_58
timestamp 1719173892
transform 1 0 -541550 0 1 -76783
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_59
timestamp 1719173892
transform 1 0 -539928 0 1 -76779
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_60
timestamp 1719173892
transform 1 0 -546066 0 1 -76783
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_61
timestamp 1719173892
transform 1 0 -544444 0 1 -76779
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_62
timestamp 1719173892
transform 1 0 -550582 0 1 -76783
box 555256 92202 556228 92502
use cv3_via2_36cut  cv3_via2_36cut_63
timestamp 1719173892
transform 1 0 -548960 0 1 -76779
box 555256 92202 556228 92502
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_0 ../ip/sky130_ef_ip__analog_switches/mag
array 0 9 -4516 0 1 4633
timestamp 1724439637
transform -1 0 3470 0 1 1481
box -4 -600 3538 3648
use simplest_analog_switch_ena1v8  simplest_analog_switch_ena1v8_1
array 0 5 -4516 0 1 4633
timestamp 1724439637
transform -1 0 3470 0 1 10747
box -4 -600 3538 3648
<< labels >>
flabel metal3 -310 15572 -310 15572 0 FreeSans 960 0 0 0 amuxbusA
flabel metal3 -260 10930 -260 10930 0 FreeSans 960 0 0 0 amuxbusB
flabel metal3 -246 6286 -246 6286 0 FreeSans 960 0 0 0 analog0
flabel metal3 -234 1674 -234 1674 0 FreeSans 960 0 0 0 analog1
flabel metal2 44342 1776 44342 1776 0 FreeSans 960 90 0 0 dac0
flabel metal2 40220 2118 40220 2118 0 FreeSans 960 90 0 0 dac1
flabel metal2 39826 2146 39826 2146 0 FreeSans 960 90 0 0 adc0
flabel metal2 35710 2188 35710 2188 0 FreeSans 960 90 0 0 adc1
flabel metal2 35298 2194 35298 2194 0 FreeSans 960 90 0 0 comp_p
flabel metal2 31178 2208 31178 2208 0 FreeSans 960 90 0 0 comp_n
flabel metal2 30786 2198 30786 2198 0 FreeSans 960 90 0 0 ulpcomp_p
flabel metal2 26674 2184 26674 2184 0 FreeSans 960 90 0 0 ulpcomp_n
flabel metal2 26272 2202 26272 2202 0 FreeSans 960 90 0 0 left_instramp_n
flabel metal2 22170 2220 22170 2220 0 FreeSans 960 90 0 0 left_instramp_p
flabel metal2 21776 2234 21776 2234 0 FreeSans 960 90 0 0 left_hgbw_opamp_n
flabel metal2 17640 2262 17640 2262 0 FreeSans 960 90 0 0 left_hgbw_opamp_p
flabel metal2 17228 2272 17228 2272 0 FreeSans 960 90 0 0 left_lp_opamp_n
flabel metal2 13132 2258 13132 2258 0 FreeSans 960 90 0 0 left_lp_opamp_p
flabel metal2 12730 2276 12730 2276 0 FreeSans 960 90 0 0 right_lp_opamp_n
flabel metal2 8616 2248 8616 2248 0 FreeSans 960 90 0 0 right_lp_opamp_p
flabel metal2 8218 2276 8218 2276 0 FreeSans 960 90 0 0 right_hgbw_opamp_n
flabel metal2 4082 2216 4082 2216 0 FreeSans 960 90 0 0 right_hgbw_opamp_p
flabel metal2 3688 2240 3688 2240 0 FreeSans 960 90 0 0 right_instramp_n
flabel metal2 -420 2618 -420 2618 0 FreeSans 960 90 0 0 right_instramp_p
flabel metal4 -650 8116 -650 8116 0 FreeSans 1600 90 0 0 vssa0
flabel metal4 3892 7804 3892 7804 0 FreeSans 1600 90 0 0 vdda0
flabel metal4 8428 7780 8428 7780 0 FreeSans 1600 90 0 0 vssd0
flabel metal4 12906 7780 12906 7780 0 FreeSans 1600 90 0 0 vccd0
<< end >>
