magic
tech sky130A
timestamp 1719106980
<< checkpaint >>
rect 284143 33430 284270 33555
<< metal2 >>
rect 284143 33550 284270 33555
rect 284143 33435 284148 33550
rect 284265 33435 284270 33550
rect 284143 33430 284270 33435
<< via2 >>
rect 284148 33435 284265 33550
<< metal3 >>
rect 284143 33550 284270 33555
rect 284143 33435 284148 33550
rect 284265 33435 284270 33550
rect 284143 33430 284270 33435
<< end >>
