magic
tech sky130A
timestamp 1723648899
<< checkpaint >>
rect 7434 10000 9142 10630
rect 0 1593 9142 10000
rect -630 874 9142 1593
rect -630 852 9183 874
rect -630 -640 9212 852
rect -630 -10630 9142 -640
<< metal4 >>
rect 0 -9779 64 10000
rect 128 -10000 192 10000
rect 256 -9779 320 10000
rect 384 -10000 448 10000
rect 512 -9779 576 10000
rect 640 -10000 704 10000
rect 768 -9779 832 10000
rect 896 -10000 960 10000
rect 1024 -9779 1088 10000
rect 1152 -10000 1216 10000
rect 1280 -9779 1344 10000
rect 1408 -10000 1472 10000
rect 1536 -9779 1600 10000
rect 1664 -10000 1728 10000
rect 1792 -9779 1856 10000
rect 1920 -10000 1984 10000
rect 2048 -9779 2112 10000
rect 2176 -10000 2240 10000
rect 2304 -9779 2368 10000
rect 2432 -10000 2496 10000
rect 2560 -9779 2624 10000
rect 2688 -10000 2752 10000
rect 2816 -9779 2880 10000
rect 2944 -10000 3008 10000
rect 3072 -9779 3136 10000
rect 3200 -10000 3264 10000
rect 3328 -9779 3392 10000
rect 3456 -10000 3520 10000
rect 3584 -9779 3648 10000
rect 3712 -10000 3776 10000
rect 3840 -9779 3904 10000
rect 3968 -10000 4032 10000
rect 4096 -9779 4160 10000
rect 4224 -10000 4288 10000
rect 4352 -9779 4416 10000
rect 4480 -10000 4544 10000
rect 4608 -9779 4672 10000
rect 4736 -10000 4800 10000
rect 4864 -9779 4928 10000
rect 4992 -10000 5056 10000
rect 5120 -9779 5184 10000
rect 5248 -10000 5312 10000
rect 5376 -9779 5440 10000
rect 5504 -10000 5568 10000
rect 5632 -9779 5696 10000
rect 5760 -10000 5824 10000
rect 5888 -9779 5952 10000
rect 6016 -10000 6080 10000
rect 6144 -9779 6208 10000
rect 6272 -10000 6336 10000
rect 6400 -9779 6464 10000
rect 6528 -10000 6592 10000
rect 6656 -9779 6720 10000
rect 6784 -10000 6848 10000
rect 6912 -9779 6976 10000
rect 7040 -10000 7104 10000
rect 7168 -9779 7232 10000
rect 7296 -10000 7360 10000
rect 7424 -9779 7488 10000
rect 7552 -10000 7616 10000
rect 7680 -9779 7744 10000
rect 7808 -10000 7872 10000
rect 7936 -9778 8000 10000
rect 8064 -10000 8128 10000
rect 8192 -9779 8256 10000
rect 8320 -10000 8384 10000
rect 8448 -9778 8512 10000
<< properties >>
string FIXED_BBOX 0 0 8000 10000
string LEFclass COVER
<< end >>
