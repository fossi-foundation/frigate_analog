magic
tech sky130A
magscale 1 2
timestamp 1717866854
<< checkpaint >>
rect -1260 -1260 242413 5558
<< metal2 >>
rect 245253 11115 245514 11136
rect 245253 10767 245278 11115
rect 245490 10767 245514 11115
rect 245253 10742 245514 10767
rect 245686 11113 245947 11135
rect 245686 10765 245714 11113
rect 245926 10765 245947 11113
rect 245686 10741 245947 10765
rect 254670 11097 254931 11119
rect 254670 10749 254695 11097
rect 254907 10749 254931 11097
rect 254670 10725 254931 10749
rect 277969 11018 278236 11042
rect 277969 10640 277993 11018
rect 278214 10640 278236 11018
rect 277969 10622 278236 10640
<< via2 >>
rect 245278 10767 245490 11115
rect 245714 10765 245926 11113
rect 254695 10749 254907 11097
rect 277993 10640 278214 11018
<< metal3 >>
rect 277861 11210 278236 11235
rect 245253 11115 245514 11136
rect 245253 10767 245278 11115
rect 245490 10767 245514 11115
rect 245253 10742 245514 10767
rect 245686 11113 245947 11135
rect 245686 10765 245714 11113
rect 245926 10765 245947 11113
rect 245686 10741 245947 10765
rect 254670 11097 254931 11119
rect 254670 10749 254695 11097
rect 254907 10749 254931 11097
rect 254670 10725 254931 10749
rect 277861 10641 277887 11210
rect 278206 11018 278236 11210
rect 277861 10640 277993 10641
rect 278214 10640 278236 11018
rect 277861 10621 278236 10640
<< via3 >>
rect 245278 10767 245490 11115
rect 245714 10765 245926 11113
rect 254695 10749 254907 11097
rect 277887 11018 278206 11210
rect 277887 10641 277993 11018
rect 277993 10641 278206 11018
<< metal4 >>
rect 238008 2797 238328 22533
rect 238662 21192 239042 21572
rect 238708 2441 239028 21192
rect 238679 2061 239059 2441
rect 239408 1431 239728 20462
rect 240078 19200 240458 19580
rect 240108 1047 240428 19200
rect 240059 667 240439 1047
rect 240808 39 241128 18624
rect 245208 17578 245564 17579
rect 245197 17198 245577 17578
rect 245241 11115 245526 17198
rect 245628 15204 246008 15584
rect 245241 10767 245278 11115
rect 245490 10767 245526 11115
rect 245241 10731 245526 10767
rect 245667 11113 245956 15204
rect 254608 13197 254988 13577
rect 245667 10765 245714 11113
rect 245926 10765 245956 11113
rect 245667 10723 245956 10765
rect 254651 11097 254951 13197
rect 277862 11569 278236 11603
rect 277858 11232 278236 11569
rect 254651 10749 254695 11097
rect 254907 10749 254951 11097
rect 254651 10708 254951 10749
rect 277862 11210 278236 11232
rect 277862 10641 277887 11210
rect 278206 10641 278236 11210
rect 277862 10622 278236 10641
<< metal5 >>
rect 238443 22235 302118 22555
rect 239042 21235 302118 21555
rect 239955 20235 302118 20555
rect 240458 19235 302118 19555
rect 240889 18235 302118 18555
rect 245577 17235 302118 17555
rect 246090 16235 302118 16555
rect 246008 15235 302118 15555
rect 246496 14235 302118 14555
rect 254988 13235 302118 13555
rect 255582 12235 302118 12555
rect 278235 11235 302118 11555
rect 278613 10235 302118 10555
rect 0 2582 238034 2902
rect 0 1940 238740 2260
rect 0 1300 239404 1620
rect 0 660 240220 980
rect 0 18 241153 338
use cv3_via4_2cut  cv3_via4_2cut_0
timestamp 1717863568
transform 1 0 277855 0 1 11205
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_1
timestamp 1717863568
transform 1 0 254608 0 1 13197
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_2
timestamp 1717863568
transform 1 0 245628 0 1 15204
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_3
timestamp 1717863568
transform 1 0 245197 0 1 17198
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_4
timestamp 1717863568
transform 1 0 239403 0 1 20215
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_5
timestamp 1717863568
transform 1 0 238662 0 1 21192
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_6
timestamp 1717863568
transform 1 0 239059 0 1 1378
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_7
timestamp 1717863568
transform 1 0 237672 0 1 2768
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_8
timestamp 1717863568
transform 1 0 240078 0 1 19200
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_9
timestamp 1717863568
transform 1 0 240809 0 1 18204
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_10
timestamp 1717863568
transform 1 0 237991 0 1 22212
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_11
timestamp 1717863568
transform 1 0 240462 0 1 0
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_12
timestamp 1717863568
transform 1 0 239744 0 1 689
box 0 0 688 368
use cv3_via4_2cut  cv3_via4_2cut_13
timestamp 1717863568
transform 1 0 238357 0 1 2067
box 0 0 688 368
<< properties >>
string FIXED_BBOX 0 0 302118 22580
string LEFclass COVER
<< end >>
